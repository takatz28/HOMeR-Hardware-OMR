/*************************************************************************
 * Module name:		tri_table
 * Input arg(s):	12-bit address
 * Output arg(s):	Triangle wave sample
 * Description:		Lookup table for triangle waveform generation
 *************************************************************************/
 
`timescale 1ns / 1ps

module tri_table (
	// port declarations
	input [11:0] tri_addr,
	output reg [15:0] tri_word
	);

	always @ (tri_addr) begin
		case (tri_addr)
			12'h000: tri_word = 16'h0000;
			12'h001: tri_word = 16'h000f;
			12'h002: tri_word = 16'h001f;
			12'h003: tri_word = 16'h002f;
			12'h004: tri_word = 16'h003f;
			12'h005: tri_word = 16'h004f;
			12'h006: tri_word = 16'h005f;
			12'h007: tri_word = 16'h006f;
			12'h008: tri_word = 16'h007f;
			12'h009: tri_word = 16'h008f;
			12'h00a: tri_word = 16'h009f;
			12'h00b: tri_word = 16'h00af;
			12'h00c: tri_word = 16'h00bf;
			12'h00d: tri_word = 16'h00cf;
			12'h00e: tri_word = 16'h00df;
			12'h00f: tri_word = 16'h00ef;
			12'h010: tri_word = 16'h00ff;
			12'h011: tri_word = 16'h010f;
			12'h012: tri_word = 16'h011f;
			12'h013: tri_word = 16'h012f;
			12'h014: tri_word = 16'h013f;
			12'h015: tri_word = 16'h014f;
			12'h016: tri_word = 16'h015f;
			12'h017: tri_word = 16'h016f;
			12'h018: tri_word = 16'h017f;
			12'h019: tri_word = 16'h018f;
			12'h01a: tri_word = 16'h019f;
			12'h01b: tri_word = 16'h01af;
			12'h01c: tri_word = 16'h01bf;
			12'h01d: tri_word = 16'h01cf;
			12'h01e: tri_word = 16'h01df;
			12'h01f: tri_word = 16'h01ef;
			12'h020: tri_word = 16'h01ff;
			12'h021: tri_word = 16'h020f;
			12'h022: tri_word = 16'h021f;
			12'h023: tri_word = 16'h022f;
			12'h024: tri_word = 16'h023f;
			12'h025: tri_word = 16'h024f;
			12'h026: tri_word = 16'h025f;
			12'h027: tri_word = 16'h026f;
			12'h028: tri_word = 16'h027f;
			12'h029: tri_word = 16'h028f;
			12'h02a: tri_word = 16'h029f;
			12'h02b: tri_word = 16'h02af;
			12'h02c: tri_word = 16'h02bf;
			12'h02d: tri_word = 16'h02cf;
			12'h02e: tri_word = 16'h02df;
			12'h02f: tri_word = 16'h02ef;
			12'h030: tri_word = 16'h02ff;
			12'h031: tri_word = 16'h030f;
			12'h032: tri_word = 16'h031f;
			12'h033: tri_word = 16'h032f;
			12'h034: tri_word = 16'h033f;
			12'h035: tri_word = 16'h034f;
			12'h036: tri_word = 16'h035f;
			12'h037: tri_word = 16'h036f;
			12'h038: tri_word = 16'h037f;
			12'h039: tri_word = 16'h038f;
			12'h03a: tri_word = 16'h039f;
			12'h03b: tri_word = 16'h03af;
			12'h03c: tri_word = 16'h03bf;
			12'h03d: tri_word = 16'h03cf;
			12'h03e: tri_word = 16'h03df;
			12'h03f: tri_word = 16'h03ef;
			12'h040: tri_word = 16'h03ff;
			12'h041: tri_word = 16'h040f;
			12'h042: tri_word = 16'h041f;
			12'h043: tri_word = 16'h042f;
			12'h044: tri_word = 16'h043f;
			12'h045: tri_word = 16'h044f;
			12'h046: tri_word = 16'h045f;
			12'h047: tri_word = 16'h046f;
			12'h048: tri_word = 16'h047f;
			12'h049: tri_word = 16'h048f;
			12'h04a: tri_word = 16'h049f;
			12'h04b: tri_word = 16'h04af;
			12'h04c: tri_word = 16'h04bf;
			12'h04d: tri_word = 16'h04cf;
			12'h04e: tri_word = 16'h04df;
			12'h04f: tri_word = 16'h04ef;
			12'h050: tri_word = 16'h04ff;
			12'h051: tri_word = 16'h050f;
			12'h052: tri_word = 16'h051f;
			12'h053: tri_word = 16'h052f;
			12'h054: tri_word = 16'h053f;
			12'h055: tri_word = 16'h054f;
			12'h056: tri_word = 16'h055f;
			12'h057: tri_word = 16'h056f;
			12'h058: tri_word = 16'h057f;
			12'h059: tri_word = 16'h058f;
			12'h05a: tri_word = 16'h059f;
			12'h05b: tri_word = 16'h05af;
			12'h05c: tri_word = 16'h05bf;
			12'h05d: tri_word = 16'h05cf;
			12'h05e: tri_word = 16'h05df;
			12'h05f: tri_word = 16'h05ef;
			12'h060: tri_word = 16'h05ff;
			12'h061: tri_word = 16'h060f;
			12'h062: tri_word = 16'h061f;
			12'h063: tri_word = 16'h062f;
			12'h064: tri_word = 16'h063f;
			12'h065: tri_word = 16'h064f;
			12'h066: tri_word = 16'h065f;
			12'h067: tri_word = 16'h066f;
			12'h068: tri_word = 16'h067f;
			12'h069: tri_word = 16'h068f;
			12'h06a: tri_word = 16'h069f;
			12'h06b: tri_word = 16'h06af;
			12'h06c: tri_word = 16'h06bf;
			12'h06d: tri_word = 16'h06cf;
			12'h06e: tri_word = 16'h06df;
			12'h06f: tri_word = 16'h06ef;
			12'h070: tri_word = 16'h06ff;
			12'h071: tri_word = 16'h070f;
			12'h072: tri_word = 16'h071f;
			12'h073: tri_word = 16'h072f;
			12'h074: tri_word = 16'h073f;
			12'h075: tri_word = 16'h074f;
			12'h076: tri_word = 16'h075f;
			12'h077: tri_word = 16'h076f;
			12'h078: tri_word = 16'h077f;
			12'h079: tri_word = 16'h078f;
			12'h07a: tri_word = 16'h079f;
			12'h07b: tri_word = 16'h07af;
			12'h07c: tri_word = 16'h07bf;
			12'h07d: tri_word = 16'h07cf;
			12'h07e: tri_word = 16'h07df;
			12'h07f: tri_word = 16'h07ef;
			12'h080: tri_word = 16'h07ff;
			12'h081: tri_word = 16'h080f;
			12'h082: tri_word = 16'h081f;
			12'h083: tri_word = 16'h082f;
			12'h084: tri_word = 16'h083f;
			12'h085: tri_word = 16'h084f;
			12'h086: tri_word = 16'h085f;
			12'h087: tri_word = 16'h086f;
			12'h088: tri_word = 16'h087f;
			12'h089: tri_word = 16'h088f;
			12'h08a: tri_word = 16'h089f;
			12'h08b: tri_word = 16'h08af;
			12'h08c: tri_word = 16'h08bf;
			12'h08d: tri_word = 16'h08cf;
			12'h08e: tri_word = 16'h08df;
			12'h08f: tri_word = 16'h08ef;
			12'h090: tri_word = 16'h08ff;
			12'h091: tri_word = 16'h090f;
			12'h092: tri_word = 16'h091f;
			12'h093: tri_word = 16'h092f;
			12'h094: tri_word = 16'h093f;
			12'h095: tri_word = 16'h094f;
			12'h096: tri_word = 16'h095f;
			12'h097: tri_word = 16'h096f;
			12'h098: tri_word = 16'h097f;
			12'h099: tri_word = 16'h098f;
			12'h09a: tri_word = 16'h099f;
			12'h09b: tri_word = 16'h09af;
			12'h09c: tri_word = 16'h09bf;
			12'h09d: tri_word = 16'h09cf;
			12'h09e: tri_word = 16'h09df;
			12'h09f: tri_word = 16'h09ef;
			12'h0a0: tri_word = 16'h09ff;
			12'h0a1: tri_word = 16'h0a0f;
			12'h0a2: tri_word = 16'h0a1f;
			12'h0a3: tri_word = 16'h0a2f;
			12'h0a4: tri_word = 16'h0a3f;
			12'h0a5: tri_word = 16'h0a4f;
			12'h0a6: tri_word = 16'h0a5f;
			12'h0a7: tri_word = 16'h0a6f;
			12'h0a8: tri_word = 16'h0a7f;
			12'h0a9: tri_word = 16'h0a8f;
			12'h0aa: tri_word = 16'h0a9f;
			12'h0ab: tri_word = 16'h0aaf;
			12'h0ac: tri_word = 16'h0abf;
			12'h0ad: tri_word = 16'h0acf;
			12'h0ae: tri_word = 16'h0adf;
			12'h0af: tri_word = 16'h0aef;
			12'h0b0: tri_word = 16'h0aff;
			12'h0b1: tri_word = 16'h0b0f;
			12'h0b2: tri_word = 16'h0b1f;
			12'h0b3: tri_word = 16'h0b2f;
			12'h0b4: tri_word = 16'h0b3f;
			12'h0b5: tri_word = 16'h0b4f;
			12'h0b6: tri_word = 16'h0b5f;
			12'h0b7: tri_word = 16'h0b6f;
			12'h0b8: tri_word = 16'h0b7f;
			12'h0b9: tri_word = 16'h0b8f;
			12'h0ba: tri_word = 16'h0b9f;
			12'h0bb: tri_word = 16'h0baf;
			12'h0bc: tri_word = 16'h0bbf;
			12'h0bd: tri_word = 16'h0bcf;
			12'h0be: tri_word = 16'h0bdf;
			12'h0bf: tri_word = 16'h0bef;
			12'h0c0: tri_word = 16'h0bff;
			12'h0c1: tri_word = 16'h0c0f;
			12'h0c2: tri_word = 16'h0c1f;
			12'h0c3: tri_word = 16'h0c2f;
			12'h0c4: tri_word = 16'h0c3f;
			12'h0c5: tri_word = 16'h0c4f;
			12'h0c6: tri_word = 16'h0c5f;
			12'h0c7: tri_word = 16'h0c6f;
			12'h0c8: tri_word = 16'h0c7f;
			12'h0c9: tri_word = 16'h0c8f;
			12'h0ca: tri_word = 16'h0c9f;
			12'h0cb: tri_word = 16'h0caf;
			12'h0cc: tri_word = 16'h0cbf;
			12'h0cd: tri_word = 16'h0ccf;
			12'h0ce: tri_word = 16'h0cdf;
			12'h0cf: tri_word = 16'h0cef;
			12'h0d0: tri_word = 16'h0cff;
			12'h0d1: tri_word = 16'h0d0f;
			12'h0d2: tri_word = 16'h0d1f;
			12'h0d3: tri_word = 16'h0d2f;
			12'h0d4: tri_word = 16'h0d3f;
			12'h0d5: tri_word = 16'h0d4f;
			12'h0d6: tri_word = 16'h0d5f;
			12'h0d7: tri_word = 16'h0d6f;
			12'h0d8: tri_word = 16'h0d7f;
			12'h0d9: tri_word = 16'h0d8f;
			12'h0da: tri_word = 16'h0d9f;
			12'h0db: tri_word = 16'h0daf;
			12'h0dc: tri_word = 16'h0dbf;
			12'h0dd: tri_word = 16'h0dcf;
			12'h0de: tri_word = 16'h0ddf;
			12'h0df: tri_word = 16'h0def;
			12'h0e0: tri_word = 16'h0dff;
			12'h0e1: tri_word = 16'h0e0f;
			12'h0e2: tri_word = 16'h0e1f;
			12'h0e3: tri_word = 16'h0e2f;
			12'h0e4: tri_word = 16'h0e3f;
			12'h0e5: tri_word = 16'h0e4f;
			12'h0e6: tri_word = 16'h0e5f;
			12'h0e7: tri_word = 16'h0e6f;
			12'h0e8: tri_word = 16'h0e7f;
			12'h0e9: tri_word = 16'h0e8f;
			12'h0ea: tri_word = 16'h0e9f;
			12'h0eb: tri_word = 16'h0eaf;
			12'h0ec: tri_word = 16'h0ebf;
			12'h0ed: tri_word = 16'h0ecf;
			12'h0ee: tri_word = 16'h0edf;
			12'h0ef: tri_word = 16'h0eef;
			12'h0f0: tri_word = 16'h0eff;
			12'h0f1: tri_word = 16'h0f0f;
			12'h0f2: tri_word = 16'h0f1f;
			12'h0f3: tri_word = 16'h0f2f;
			12'h0f4: tri_word = 16'h0f3f;
			12'h0f5: tri_word = 16'h0f4f;
			12'h0f6: tri_word = 16'h0f5f;
			12'h0f7: tri_word = 16'h0f6f;
			12'h0f8: tri_word = 16'h0f7f;
			12'h0f9: tri_word = 16'h0f8f;
			12'h0fa: tri_word = 16'h0f9f;
			12'h0fb: tri_word = 16'h0faf;
			12'h0fc: tri_word = 16'h0fbf;
			12'h0fd: tri_word = 16'h0fcf;
			12'h0fe: tri_word = 16'h0fdf;
			12'h0ff: tri_word = 16'h0fef;
			12'h100: tri_word = 16'h0fff;
			12'h101: tri_word = 16'h100f;
			12'h102: tri_word = 16'h101f;
			12'h103: tri_word = 16'h102f;
			12'h104: tri_word = 16'h103f;
			12'h105: tri_word = 16'h104f;
			12'h106: tri_word = 16'h105f;
			12'h107: tri_word = 16'h106f;
			12'h108: tri_word = 16'h107f;
			12'h109: tri_word = 16'h108f;
			12'h10a: tri_word = 16'h109f;
			12'h10b: tri_word = 16'h10af;
			12'h10c: tri_word = 16'h10bf;
			12'h10d: tri_word = 16'h10cf;
			12'h10e: tri_word = 16'h10df;
			12'h10f: tri_word = 16'h10ef;
			12'h110: tri_word = 16'h10ff;
			12'h111: tri_word = 16'h110f;
			12'h112: tri_word = 16'h111f;
			12'h113: tri_word = 16'h112f;
			12'h114: tri_word = 16'h113f;
			12'h115: tri_word = 16'h114f;
			12'h116: tri_word = 16'h115f;
			12'h117: tri_word = 16'h116f;
			12'h118: tri_word = 16'h117f;
			12'h119: tri_word = 16'h118f;
			12'h11a: tri_word = 16'h119f;
			12'h11b: tri_word = 16'h11af;
			12'h11c: tri_word = 16'h11bf;
			12'h11d: tri_word = 16'h11cf;
			12'h11e: tri_word = 16'h11df;
			12'h11f: tri_word = 16'h11ef;
			12'h120: tri_word = 16'h11ff;
			12'h121: tri_word = 16'h120f;
			12'h122: tri_word = 16'h121f;
			12'h123: tri_word = 16'h122f;
			12'h124: tri_word = 16'h123f;
			12'h125: tri_word = 16'h124f;
			12'h126: tri_word = 16'h125f;
			12'h127: tri_word = 16'h126f;
			12'h128: tri_word = 16'h127f;
			12'h129: tri_word = 16'h128f;
			12'h12a: tri_word = 16'h129f;
			12'h12b: tri_word = 16'h12af;
			12'h12c: tri_word = 16'h12bf;
			12'h12d: tri_word = 16'h12cf;
			12'h12e: tri_word = 16'h12df;
			12'h12f: tri_word = 16'h12ef;
			12'h130: tri_word = 16'h12ff;
			12'h131: tri_word = 16'h130f;
			12'h132: tri_word = 16'h131f;
			12'h133: tri_word = 16'h132f;
			12'h134: tri_word = 16'h133f;
			12'h135: tri_word = 16'h134f;
			12'h136: tri_word = 16'h135f;
			12'h137: tri_word = 16'h136f;
			12'h138: tri_word = 16'h137f;
			12'h139: tri_word = 16'h138f;
			12'h13a: tri_word = 16'h139f;
			12'h13b: tri_word = 16'h13af;
			12'h13c: tri_word = 16'h13bf;
			12'h13d: tri_word = 16'h13cf;
			12'h13e: tri_word = 16'h13df;
			12'h13f: tri_word = 16'h13ef;
			12'h140: tri_word = 16'h13ff;
			12'h141: tri_word = 16'h140f;
			12'h142: tri_word = 16'h141f;
			12'h143: tri_word = 16'h142f;
			12'h144: tri_word = 16'h143f;
			12'h145: tri_word = 16'h144f;
			12'h146: tri_word = 16'h145f;
			12'h147: tri_word = 16'h146f;
			12'h148: tri_word = 16'h147f;
			12'h149: tri_word = 16'h148f;
			12'h14a: tri_word = 16'h149f;
			12'h14b: tri_word = 16'h14af;
			12'h14c: tri_word = 16'h14bf;
			12'h14d: tri_word = 16'h14cf;
			12'h14e: tri_word = 16'h14df;
			12'h14f: tri_word = 16'h14ef;
			12'h150: tri_word = 16'h14ff;
			12'h151: tri_word = 16'h150f;
			12'h152: tri_word = 16'h151f;
			12'h153: tri_word = 16'h152f;
			12'h154: tri_word = 16'h153f;
			12'h155: tri_word = 16'h154f;
			12'h156: tri_word = 16'h155f;
			12'h157: tri_word = 16'h156f;
			12'h158: tri_word = 16'h157f;
			12'h159: tri_word = 16'h158f;
			12'h15a: tri_word = 16'h159f;
			12'h15b: tri_word = 16'h15af;
			12'h15c: tri_word = 16'h15bf;
			12'h15d: tri_word = 16'h15cf;
			12'h15e: tri_word = 16'h15df;
			12'h15f: tri_word = 16'h15ef;
			12'h160: tri_word = 16'h15ff;
			12'h161: tri_word = 16'h160f;
			12'h162: tri_word = 16'h161f;
			12'h163: tri_word = 16'h162f;
			12'h164: tri_word = 16'h163f;
			12'h165: tri_word = 16'h164f;
			12'h166: tri_word = 16'h165f;
			12'h167: tri_word = 16'h166f;
			12'h168: tri_word = 16'h167f;
			12'h169: tri_word = 16'h168f;
			12'h16a: tri_word = 16'h169f;
			12'h16b: tri_word = 16'h16af;
			12'h16c: tri_word = 16'h16bf;
			12'h16d: tri_word = 16'h16cf;
			12'h16e: tri_word = 16'h16df;
			12'h16f: tri_word = 16'h16ef;
			12'h170: tri_word = 16'h16ff;
			12'h171: tri_word = 16'h170f;
			12'h172: tri_word = 16'h171f;
			12'h173: tri_word = 16'h172f;
			12'h174: tri_word = 16'h173f;
			12'h175: tri_word = 16'h174f;
			12'h176: tri_word = 16'h175f;
			12'h177: tri_word = 16'h176f;
			12'h178: tri_word = 16'h177f;
			12'h179: tri_word = 16'h178f;
			12'h17a: tri_word = 16'h179f;
			12'h17b: tri_word = 16'h17af;
			12'h17c: tri_word = 16'h17bf;
			12'h17d: tri_word = 16'h17cf;
			12'h17e: tri_word = 16'h17df;
			12'h17f: tri_word = 16'h17ef;
			12'h180: tri_word = 16'h17ff;
			12'h181: tri_word = 16'h180f;
			12'h182: tri_word = 16'h181f;
			12'h183: tri_word = 16'h182f;
			12'h184: tri_word = 16'h183f;
			12'h185: tri_word = 16'h184f;
			12'h186: tri_word = 16'h185f;
			12'h187: tri_word = 16'h186f;
			12'h188: tri_word = 16'h187f;
			12'h189: tri_word = 16'h188f;
			12'h18a: tri_word = 16'h189f;
			12'h18b: tri_word = 16'h18af;
			12'h18c: tri_word = 16'h18bf;
			12'h18d: tri_word = 16'h18cf;
			12'h18e: tri_word = 16'h18df;
			12'h18f: tri_word = 16'h18ef;
			12'h190: tri_word = 16'h18ff;
			12'h191: tri_word = 16'h190f;
			12'h192: tri_word = 16'h191f;
			12'h193: tri_word = 16'h192f;
			12'h194: tri_word = 16'h193f;
			12'h195: tri_word = 16'h194f;
			12'h196: tri_word = 16'h195f;
			12'h197: tri_word = 16'h196f;
			12'h198: tri_word = 16'h197f;
			12'h199: tri_word = 16'h198f;
			12'h19a: tri_word = 16'h199f;
			12'h19b: tri_word = 16'h19af;
			12'h19c: tri_word = 16'h19bf;
			12'h19d: tri_word = 16'h19cf;
			12'h19e: tri_word = 16'h19df;
			12'h19f: tri_word = 16'h19ef;
			12'h1a0: tri_word = 16'h19ff;
			12'h1a1: tri_word = 16'h1a0f;
			12'h1a2: tri_word = 16'h1a1f;
			12'h1a3: tri_word = 16'h1a2f;
			12'h1a4: tri_word = 16'h1a3f;
			12'h1a5: tri_word = 16'h1a4f;
			12'h1a6: tri_word = 16'h1a5f;
			12'h1a7: tri_word = 16'h1a6f;
			12'h1a8: tri_word = 16'h1a7f;
			12'h1a9: tri_word = 16'h1a8f;
			12'h1aa: tri_word = 16'h1a9f;
			12'h1ab: tri_word = 16'h1aaf;
			12'h1ac: tri_word = 16'h1abf;
			12'h1ad: tri_word = 16'h1acf;
			12'h1ae: tri_word = 16'h1adf;
			12'h1af: tri_word = 16'h1aef;
			12'h1b0: tri_word = 16'h1aff;
			12'h1b1: tri_word = 16'h1b0f;
			12'h1b2: tri_word = 16'h1b1f;
			12'h1b3: tri_word = 16'h1b2f;
			12'h1b4: tri_word = 16'h1b3f;
			12'h1b5: tri_word = 16'h1b4f;
			12'h1b6: tri_word = 16'h1b5f;
			12'h1b7: tri_word = 16'h1b6f;
			12'h1b8: tri_word = 16'h1b7f;
			12'h1b9: tri_word = 16'h1b8f;
			12'h1ba: tri_word = 16'h1b9f;
			12'h1bb: tri_word = 16'h1baf;
			12'h1bc: tri_word = 16'h1bbf;
			12'h1bd: tri_word = 16'h1bcf;
			12'h1be: tri_word = 16'h1bdf;
			12'h1bf: tri_word = 16'h1bef;
			12'h1c0: tri_word = 16'h1bff;
			12'h1c1: tri_word = 16'h1c0f;
			12'h1c2: tri_word = 16'h1c1f;
			12'h1c3: tri_word = 16'h1c2f;
			12'h1c4: tri_word = 16'h1c3f;
			12'h1c5: tri_word = 16'h1c4f;
			12'h1c6: tri_word = 16'h1c5f;
			12'h1c7: tri_word = 16'h1c6f;
			12'h1c8: tri_word = 16'h1c7f;
			12'h1c9: tri_word = 16'h1c8f;
			12'h1ca: tri_word = 16'h1c9f;
			12'h1cb: tri_word = 16'h1caf;
			12'h1cc: tri_word = 16'h1cbf;
			12'h1cd: tri_word = 16'h1ccf;
			12'h1ce: tri_word = 16'h1cdf;
			12'h1cf: tri_word = 16'h1cef;
			12'h1d0: tri_word = 16'h1cff;
			12'h1d1: tri_word = 16'h1d0f;
			12'h1d2: tri_word = 16'h1d1f;
			12'h1d3: tri_word = 16'h1d2f;
			12'h1d4: tri_word = 16'h1d3f;
			12'h1d5: tri_word = 16'h1d4f;
			12'h1d6: tri_word = 16'h1d5f;
			12'h1d7: tri_word = 16'h1d6f;
			12'h1d8: tri_word = 16'h1d7f;
			12'h1d9: tri_word = 16'h1d8f;
			12'h1da: tri_word = 16'h1d9f;
			12'h1db: tri_word = 16'h1daf;
			12'h1dc: tri_word = 16'h1dbf;
			12'h1dd: tri_word = 16'h1dcf;
			12'h1de: tri_word = 16'h1ddf;
			12'h1df: tri_word = 16'h1def;
			12'h1e0: tri_word = 16'h1dff;
			12'h1e1: tri_word = 16'h1e0f;
			12'h1e2: tri_word = 16'h1e1f;
			12'h1e3: tri_word = 16'h1e2f;
			12'h1e4: tri_word = 16'h1e3f;
			12'h1e5: tri_word = 16'h1e4f;
			12'h1e6: tri_word = 16'h1e5f;
			12'h1e7: tri_word = 16'h1e6f;
			12'h1e8: tri_word = 16'h1e7f;
			12'h1e9: tri_word = 16'h1e8f;
			12'h1ea: tri_word = 16'h1e9f;
			12'h1eb: tri_word = 16'h1eaf;
			12'h1ec: tri_word = 16'h1ebf;
			12'h1ed: tri_word = 16'h1ecf;
			12'h1ee: tri_word = 16'h1edf;
			12'h1ef: tri_word = 16'h1eef;
			12'h1f0: tri_word = 16'h1eff;
			12'h1f1: tri_word = 16'h1f0f;
			12'h1f2: tri_word = 16'h1f1f;
			12'h1f3: tri_word = 16'h1f2f;
			12'h1f4: tri_word = 16'h1f3f;
			12'h1f5: tri_word = 16'h1f4f;
			12'h1f6: tri_word = 16'h1f5f;
			12'h1f7: tri_word = 16'h1f6f;
			12'h1f8: tri_word = 16'h1f7f;
			12'h1f9: tri_word = 16'h1f8f;
			12'h1fa: tri_word = 16'h1f9f;
			12'h1fb: tri_word = 16'h1faf;
			12'h1fc: tri_word = 16'h1fbf;
			12'h1fd: tri_word = 16'h1fcf;
			12'h1fe: tri_word = 16'h1fdf;
			12'h1ff: tri_word = 16'h1fef;
			12'h200: tri_word = 16'h1fff;
			12'h201: tri_word = 16'h200f;
			12'h202: tri_word = 16'h201f;
			12'h203: tri_word = 16'h202f;
			12'h204: tri_word = 16'h203f;
			12'h205: tri_word = 16'h204f;
			12'h206: tri_word = 16'h205f;
			12'h207: tri_word = 16'h206f;
			12'h208: tri_word = 16'h207f;
			12'h209: tri_word = 16'h208f;
			12'h20a: tri_word = 16'h209f;
			12'h20b: tri_word = 16'h20af;
			12'h20c: tri_word = 16'h20bf;
			12'h20d: tri_word = 16'h20cf;
			12'h20e: tri_word = 16'h20df;
			12'h20f: tri_word = 16'h20ef;
			12'h210: tri_word = 16'h20ff;
			12'h211: tri_word = 16'h210f;
			12'h212: tri_word = 16'h211f;
			12'h213: tri_word = 16'h212f;
			12'h214: tri_word = 16'h213f;
			12'h215: tri_word = 16'h214f;
			12'h216: tri_word = 16'h215f;
			12'h217: tri_word = 16'h216f;
			12'h218: tri_word = 16'h217f;
			12'h219: tri_word = 16'h218f;
			12'h21a: tri_word = 16'h219f;
			12'h21b: tri_word = 16'h21af;
			12'h21c: tri_word = 16'h21bf;
			12'h21d: tri_word = 16'h21cf;
			12'h21e: tri_word = 16'h21df;
			12'h21f: tri_word = 16'h21ef;
			12'h220: tri_word = 16'h21ff;
			12'h221: tri_word = 16'h220f;
			12'h222: tri_word = 16'h221f;
			12'h223: tri_word = 16'h222f;
			12'h224: tri_word = 16'h223f;
			12'h225: tri_word = 16'h224f;
			12'h226: tri_word = 16'h225f;
			12'h227: tri_word = 16'h226f;
			12'h228: tri_word = 16'h227f;
			12'h229: tri_word = 16'h228f;
			12'h22a: tri_word = 16'h229f;
			12'h22b: tri_word = 16'h22af;
			12'h22c: tri_word = 16'h22bf;
			12'h22d: tri_word = 16'h22cf;
			12'h22e: tri_word = 16'h22df;
			12'h22f: tri_word = 16'h22ef;
			12'h230: tri_word = 16'h22ff;
			12'h231: tri_word = 16'h230f;
			12'h232: tri_word = 16'h231f;
			12'h233: tri_word = 16'h232f;
			12'h234: tri_word = 16'h233f;
			12'h235: tri_word = 16'h234f;
			12'h236: tri_word = 16'h235f;
			12'h237: tri_word = 16'h236f;
			12'h238: tri_word = 16'h237f;
			12'h239: tri_word = 16'h238f;
			12'h23a: tri_word = 16'h239f;
			12'h23b: tri_word = 16'h23af;
			12'h23c: tri_word = 16'h23bf;
			12'h23d: tri_word = 16'h23cf;
			12'h23e: tri_word = 16'h23df;
			12'h23f: tri_word = 16'h23ef;
			12'h240: tri_word = 16'h23ff;
			12'h241: tri_word = 16'h240f;
			12'h242: tri_word = 16'h241f;
			12'h243: tri_word = 16'h242f;
			12'h244: tri_word = 16'h243f;
			12'h245: tri_word = 16'h244f;
			12'h246: tri_word = 16'h245f;
			12'h247: tri_word = 16'h246f;
			12'h248: tri_word = 16'h247f;
			12'h249: tri_word = 16'h248f;
			12'h24a: tri_word = 16'h249f;
			12'h24b: tri_word = 16'h24af;
			12'h24c: tri_word = 16'h24bf;
			12'h24d: tri_word = 16'h24cf;
			12'h24e: tri_word = 16'h24df;
			12'h24f: tri_word = 16'h24ef;
			12'h250: tri_word = 16'h24ff;
			12'h251: tri_word = 16'h250f;
			12'h252: tri_word = 16'h251f;
			12'h253: tri_word = 16'h252f;
			12'h254: tri_word = 16'h253f;
			12'h255: tri_word = 16'h254f;
			12'h256: tri_word = 16'h255f;
			12'h257: tri_word = 16'h256f;
			12'h258: tri_word = 16'h257f;
			12'h259: tri_word = 16'h258f;
			12'h25a: tri_word = 16'h259f;
			12'h25b: tri_word = 16'h25af;
			12'h25c: tri_word = 16'h25bf;
			12'h25d: tri_word = 16'h25cf;
			12'h25e: tri_word = 16'h25df;
			12'h25f: tri_word = 16'h25ef;
			12'h260: tri_word = 16'h25ff;
			12'h261: tri_word = 16'h260f;
			12'h262: tri_word = 16'h261f;
			12'h263: tri_word = 16'h262f;
			12'h264: tri_word = 16'h263f;
			12'h265: tri_word = 16'h264f;
			12'h266: tri_word = 16'h265f;
			12'h267: tri_word = 16'h266f;
			12'h268: tri_word = 16'h267f;
			12'h269: tri_word = 16'h268f;
			12'h26a: tri_word = 16'h269f;
			12'h26b: tri_word = 16'h26af;
			12'h26c: tri_word = 16'h26bf;
			12'h26d: tri_word = 16'h26cf;
			12'h26e: tri_word = 16'h26df;
			12'h26f: tri_word = 16'h26ef;
			12'h270: tri_word = 16'h26ff;
			12'h271: tri_word = 16'h270f;
			12'h272: tri_word = 16'h271f;
			12'h273: tri_word = 16'h272f;
			12'h274: tri_word = 16'h273f;
			12'h275: tri_word = 16'h274f;
			12'h276: tri_word = 16'h275f;
			12'h277: tri_word = 16'h276f;
			12'h278: tri_word = 16'h277f;
			12'h279: tri_word = 16'h278f;
			12'h27a: tri_word = 16'h279f;
			12'h27b: tri_word = 16'h27af;
			12'h27c: tri_word = 16'h27bf;
			12'h27d: tri_word = 16'h27cf;
			12'h27e: tri_word = 16'h27df;
			12'h27f: tri_word = 16'h27ef;
			12'h280: tri_word = 16'h27ff;
			12'h281: tri_word = 16'h280f;
			12'h282: tri_word = 16'h281f;
			12'h283: tri_word = 16'h282f;
			12'h284: tri_word = 16'h283f;
			12'h285: tri_word = 16'h284f;
			12'h286: tri_word = 16'h285f;
			12'h287: tri_word = 16'h286f;
			12'h288: tri_word = 16'h287f;
			12'h289: tri_word = 16'h288f;
			12'h28a: tri_word = 16'h289f;
			12'h28b: tri_word = 16'h28af;
			12'h28c: tri_word = 16'h28bf;
			12'h28d: tri_word = 16'h28cf;
			12'h28e: tri_word = 16'h28df;
			12'h28f: tri_word = 16'h28ef;
			12'h290: tri_word = 16'h28ff;
			12'h291: tri_word = 16'h290f;
			12'h292: tri_word = 16'h291f;
			12'h293: tri_word = 16'h292f;
			12'h294: tri_word = 16'h293f;
			12'h295: tri_word = 16'h294f;
			12'h296: tri_word = 16'h295f;
			12'h297: tri_word = 16'h296f;
			12'h298: tri_word = 16'h297f;
			12'h299: tri_word = 16'h298f;
			12'h29a: tri_word = 16'h299f;
			12'h29b: tri_word = 16'h29af;
			12'h29c: tri_word = 16'h29bf;
			12'h29d: tri_word = 16'h29cf;
			12'h29e: tri_word = 16'h29df;
			12'h29f: tri_word = 16'h29ef;
			12'h2a0: tri_word = 16'h29ff;
			12'h2a1: tri_word = 16'h2a0f;
			12'h2a2: tri_word = 16'h2a1f;
			12'h2a3: tri_word = 16'h2a2f;
			12'h2a4: tri_word = 16'h2a3f;
			12'h2a5: tri_word = 16'h2a4f;
			12'h2a6: tri_word = 16'h2a5f;
			12'h2a7: tri_word = 16'h2a6f;
			12'h2a8: tri_word = 16'h2a7f;
			12'h2a9: tri_word = 16'h2a8f;
			12'h2aa: tri_word = 16'h2a9f;
			12'h2ab: tri_word = 16'h2aaf;
			12'h2ac: tri_word = 16'h2abf;
			12'h2ad: tri_word = 16'h2acf;
			12'h2ae: tri_word = 16'h2adf;
			12'h2af: tri_word = 16'h2aef;
			12'h2b0: tri_word = 16'h2aff;
			12'h2b1: tri_word = 16'h2b0f;
			12'h2b2: tri_word = 16'h2b1f;
			12'h2b3: tri_word = 16'h2b2f;
			12'h2b4: tri_word = 16'h2b3f;
			12'h2b5: tri_word = 16'h2b4f;
			12'h2b6: tri_word = 16'h2b5f;
			12'h2b7: tri_word = 16'h2b6f;
			12'h2b8: tri_word = 16'h2b7f;
			12'h2b9: tri_word = 16'h2b8f;
			12'h2ba: tri_word = 16'h2b9f;
			12'h2bb: tri_word = 16'h2baf;
			12'h2bc: tri_word = 16'h2bbf;
			12'h2bd: tri_word = 16'h2bcf;
			12'h2be: tri_word = 16'h2bdf;
			12'h2bf: tri_word = 16'h2bef;
			12'h2c0: tri_word = 16'h2bff;
			12'h2c1: tri_word = 16'h2c0f;
			12'h2c2: tri_word = 16'h2c1f;
			12'h2c3: tri_word = 16'h2c2f;
			12'h2c4: tri_word = 16'h2c3f;
			12'h2c5: tri_word = 16'h2c4f;
			12'h2c6: tri_word = 16'h2c5f;
			12'h2c7: tri_word = 16'h2c6f;
			12'h2c8: tri_word = 16'h2c7f;
			12'h2c9: tri_word = 16'h2c8f;
			12'h2ca: tri_word = 16'h2c9f;
			12'h2cb: tri_word = 16'h2caf;
			12'h2cc: tri_word = 16'h2cbf;
			12'h2cd: tri_word = 16'h2ccf;
			12'h2ce: tri_word = 16'h2cdf;
			12'h2cf: tri_word = 16'h2cef;
			12'h2d0: tri_word = 16'h2cff;
			12'h2d1: tri_word = 16'h2d0f;
			12'h2d2: tri_word = 16'h2d1f;
			12'h2d3: tri_word = 16'h2d2f;
			12'h2d4: tri_word = 16'h2d3f;
			12'h2d5: tri_word = 16'h2d4f;
			12'h2d6: tri_word = 16'h2d5f;
			12'h2d7: tri_word = 16'h2d6f;
			12'h2d8: tri_word = 16'h2d7f;
			12'h2d9: tri_word = 16'h2d8f;
			12'h2da: tri_word = 16'h2d9f;
			12'h2db: tri_word = 16'h2daf;
			12'h2dc: tri_word = 16'h2dbf;
			12'h2dd: tri_word = 16'h2dcf;
			12'h2de: tri_word = 16'h2ddf;
			12'h2df: tri_word = 16'h2def;
			12'h2e0: tri_word = 16'h2dff;
			12'h2e1: tri_word = 16'h2e0f;
			12'h2e2: tri_word = 16'h2e1f;
			12'h2e3: tri_word = 16'h2e2f;
			12'h2e4: tri_word = 16'h2e3f;
			12'h2e5: tri_word = 16'h2e4f;
			12'h2e6: tri_word = 16'h2e5f;
			12'h2e7: tri_word = 16'h2e6f;
			12'h2e8: tri_word = 16'h2e7f;
			12'h2e9: tri_word = 16'h2e8f;
			12'h2ea: tri_word = 16'h2e9f;
			12'h2eb: tri_word = 16'h2eaf;
			12'h2ec: tri_word = 16'h2ebf;
			12'h2ed: tri_word = 16'h2ecf;
			12'h2ee: tri_word = 16'h2edf;
			12'h2ef: tri_word = 16'h2eef;
			12'h2f0: tri_word = 16'h2eff;
			12'h2f1: tri_word = 16'h2f0f;
			12'h2f2: tri_word = 16'h2f1f;
			12'h2f3: tri_word = 16'h2f2f;
			12'h2f4: tri_word = 16'h2f3f;
			12'h2f5: tri_word = 16'h2f4f;
			12'h2f6: tri_word = 16'h2f5f;
			12'h2f7: tri_word = 16'h2f6f;
			12'h2f8: tri_word = 16'h2f7f;
			12'h2f9: tri_word = 16'h2f8f;
			12'h2fa: tri_word = 16'h2f9f;
			12'h2fb: tri_word = 16'h2faf;
			12'h2fc: tri_word = 16'h2fbf;
			12'h2fd: tri_word = 16'h2fcf;
			12'h2fe: tri_word = 16'h2fdf;
			12'h2ff: tri_word = 16'h2fef;
			12'h300: tri_word = 16'h2fff;
			12'h301: tri_word = 16'h300f;
			12'h302: tri_word = 16'h301f;
			12'h303: tri_word = 16'h302f;
			12'h304: tri_word = 16'h303f;
			12'h305: tri_word = 16'h304f;
			12'h306: tri_word = 16'h305f;
			12'h307: tri_word = 16'h306f;
			12'h308: tri_word = 16'h307f;
			12'h309: tri_word = 16'h308f;
			12'h30a: tri_word = 16'h309f;
			12'h30b: tri_word = 16'h30af;
			12'h30c: tri_word = 16'h30bf;
			12'h30d: tri_word = 16'h30cf;
			12'h30e: tri_word = 16'h30df;
			12'h30f: tri_word = 16'h30ef;
			12'h310: tri_word = 16'h30ff;
			12'h311: tri_word = 16'h310f;
			12'h312: tri_word = 16'h311f;
			12'h313: tri_word = 16'h312f;
			12'h314: tri_word = 16'h313f;
			12'h315: tri_word = 16'h314f;
			12'h316: tri_word = 16'h315f;
			12'h317: tri_word = 16'h316f;
			12'h318: tri_word = 16'h317f;
			12'h319: tri_word = 16'h318f;
			12'h31a: tri_word = 16'h319f;
			12'h31b: tri_word = 16'h31af;
			12'h31c: tri_word = 16'h31bf;
			12'h31d: tri_word = 16'h31cf;
			12'h31e: tri_word = 16'h31df;
			12'h31f: tri_word = 16'h31ef;
			12'h320: tri_word = 16'h31ff;
			12'h321: tri_word = 16'h320f;
			12'h322: tri_word = 16'h321f;
			12'h323: tri_word = 16'h322f;
			12'h324: tri_word = 16'h323f;
			12'h325: tri_word = 16'h324f;
			12'h326: tri_word = 16'h325f;
			12'h327: tri_word = 16'h326f;
			12'h328: tri_word = 16'h327f;
			12'h329: tri_word = 16'h328f;
			12'h32a: tri_word = 16'h329f;
			12'h32b: tri_word = 16'h32af;
			12'h32c: tri_word = 16'h32bf;
			12'h32d: tri_word = 16'h32cf;
			12'h32e: tri_word = 16'h32df;
			12'h32f: tri_word = 16'h32ef;
			12'h330: tri_word = 16'h32ff;
			12'h331: tri_word = 16'h330f;
			12'h332: tri_word = 16'h331f;
			12'h333: tri_word = 16'h332f;
			12'h334: tri_word = 16'h333f;
			12'h335: tri_word = 16'h334f;
			12'h336: tri_word = 16'h335f;
			12'h337: tri_word = 16'h336f;
			12'h338: tri_word = 16'h337f;
			12'h339: tri_word = 16'h338f;
			12'h33a: tri_word = 16'h339f;
			12'h33b: tri_word = 16'h33af;
			12'h33c: tri_word = 16'h33bf;
			12'h33d: tri_word = 16'h33cf;
			12'h33e: tri_word = 16'h33df;
			12'h33f: tri_word = 16'h33ef;
			12'h340: tri_word = 16'h33ff;
			12'h341: tri_word = 16'h340f;
			12'h342: tri_word = 16'h341f;
			12'h343: tri_word = 16'h342f;
			12'h344: tri_word = 16'h343f;
			12'h345: tri_word = 16'h344f;
			12'h346: tri_word = 16'h345f;
			12'h347: tri_word = 16'h346f;
			12'h348: tri_word = 16'h347f;
			12'h349: tri_word = 16'h348f;
			12'h34a: tri_word = 16'h349f;
			12'h34b: tri_word = 16'h34af;
			12'h34c: tri_word = 16'h34bf;
			12'h34d: tri_word = 16'h34cf;
			12'h34e: tri_word = 16'h34df;
			12'h34f: tri_word = 16'h34ef;
			12'h350: tri_word = 16'h34ff;
			12'h351: tri_word = 16'h350f;
			12'h352: tri_word = 16'h351f;
			12'h353: tri_word = 16'h352f;
			12'h354: tri_word = 16'h353f;
			12'h355: tri_word = 16'h354f;
			12'h356: tri_word = 16'h355f;
			12'h357: tri_word = 16'h356f;
			12'h358: tri_word = 16'h357f;
			12'h359: tri_word = 16'h358f;
			12'h35a: tri_word = 16'h359f;
			12'h35b: tri_word = 16'h35af;
			12'h35c: tri_word = 16'h35bf;
			12'h35d: tri_word = 16'h35cf;
			12'h35e: tri_word = 16'h35df;
			12'h35f: tri_word = 16'h35ef;
			12'h360: tri_word = 16'h35ff;
			12'h361: tri_word = 16'h360f;
			12'h362: tri_word = 16'h361f;
			12'h363: tri_word = 16'h362f;
			12'h364: tri_word = 16'h363f;
			12'h365: tri_word = 16'h364f;
			12'h366: tri_word = 16'h365f;
			12'h367: tri_word = 16'h366f;
			12'h368: tri_word = 16'h367f;
			12'h369: tri_word = 16'h368f;
			12'h36a: tri_word = 16'h369f;
			12'h36b: tri_word = 16'h36af;
			12'h36c: tri_word = 16'h36bf;
			12'h36d: tri_word = 16'h36cf;
			12'h36e: tri_word = 16'h36df;
			12'h36f: tri_word = 16'h36ef;
			12'h370: tri_word = 16'h36ff;
			12'h371: tri_word = 16'h370f;
			12'h372: tri_word = 16'h371f;
			12'h373: tri_word = 16'h372f;
			12'h374: tri_word = 16'h373f;
			12'h375: tri_word = 16'h374f;
			12'h376: tri_word = 16'h375f;
			12'h377: tri_word = 16'h376f;
			12'h378: tri_word = 16'h377f;
			12'h379: tri_word = 16'h378f;
			12'h37a: tri_word = 16'h379f;
			12'h37b: tri_word = 16'h37af;
			12'h37c: tri_word = 16'h37bf;
			12'h37d: tri_word = 16'h37cf;
			12'h37e: tri_word = 16'h37df;
			12'h37f: tri_word = 16'h37ef;
			12'h380: tri_word = 16'h37ff;
			12'h381: tri_word = 16'h380f;
			12'h382: tri_word = 16'h381f;
			12'h383: tri_word = 16'h382f;
			12'h384: tri_word = 16'h383f;
			12'h385: tri_word = 16'h384f;
			12'h386: tri_word = 16'h385f;
			12'h387: tri_word = 16'h386f;
			12'h388: tri_word = 16'h387f;
			12'h389: tri_word = 16'h388f;
			12'h38a: tri_word = 16'h389f;
			12'h38b: tri_word = 16'h38af;
			12'h38c: tri_word = 16'h38bf;
			12'h38d: tri_word = 16'h38cf;
			12'h38e: tri_word = 16'h38df;
			12'h38f: tri_word = 16'h38ef;
			12'h390: tri_word = 16'h38ff;
			12'h391: tri_word = 16'h390f;
			12'h392: tri_word = 16'h391f;
			12'h393: tri_word = 16'h392f;
			12'h394: tri_word = 16'h393f;
			12'h395: tri_word = 16'h394f;
			12'h396: tri_word = 16'h395f;
			12'h397: tri_word = 16'h396f;
			12'h398: tri_word = 16'h397f;
			12'h399: tri_word = 16'h398f;
			12'h39a: tri_word = 16'h399f;
			12'h39b: tri_word = 16'h39af;
			12'h39c: tri_word = 16'h39bf;
			12'h39d: tri_word = 16'h39cf;
			12'h39e: tri_word = 16'h39df;
			12'h39f: tri_word = 16'h39ef;
			12'h3a0: tri_word = 16'h39ff;
			12'h3a1: tri_word = 16'h3a0f;
			12'h3a2: tri_word = 16'h3a1f;
			12'h3a3: tri_word = 16'h3a2f;
			12'h3a4: tri_word = 16'h3a3f;
			12'h3a5: tri_word = 16'h3a4f;
			12'h3a6: tri_word = 16'h3a5f;
			12'h3a7: tri_word = 16'h3a6f;
			12'h3a8: tri_word = 16'h3a7f;
			12'h3a9: tri_word = 16'h3a8f;
			12'h3aa: tri_word = 16'h3a9f;
			12'h3ab: tri_word = 16'h3aaf;
			12'h3ac: tri_word = 16'h3abf;
			12'h3ad: tri_word = 16'h3acf;
			12'h3ae: tri_word = 16'h3adf;
			12'h3af: tri_word = 16'h3aef;
			12'h3b0: tri_word = 16'h3aff;
			12'h3b1: tri_word = 16'h3b0f;
			12'h3b2: tri_word = 16'h3b1f;
			12'h3b3: tri_word = 16'h3b2f;
			12'h3b4: tri_word = 16'h3b3f;
			12'h3b5: tri_word = 16'h3b4f;
			12'h3b6: tri_word = 16'h3b5f;
			12'h3b7: tri_word = 16'h3b6f;
			12'h3b8: tri_word = 16'h3b7f;
			12'h3b9: tri_word = 16'h3b8f;
			12'h3ba: tri_word = 16'h3b9f;
			12'h3bb: tri_word = 16'h3baf;
			12'h3bc: tri_word = 16'h3bbf;
			12'h3bd: tri_word = 16'h3bcf;
			12'h3be: tri_word = 16'h3bdf;
			12'h3bf: tri_word = 16'h3bef;
			12'h3c0: tri_word = 16'h3bff;
			12'h3c1: tri_word = 16'h3c0f;
			12'h3c2: tri_word = 16'h3c1f;
			12'h3c3: tri_word = 16'h3c2f;
			12'h3c4: tri_word = 16'h3c3f;
			12'h3c5: tri_word = 16'h3c4f;
			12'h3c6: tri_word = 16'h3c5f;
			12'h3c7: tri_word = 16'h3c6f;
			12'h3c8: tri_word = 16'h3c7f;
			12'h3c9: tri_word = 16'h3c8f;
			12'h3ca: tri_word = 16'h3c9f;
			12'h3cb: tri_word = 16'h3caf;
			12'h3cc: tri_word = 16'h3cbf;
			12'h3cd: tri_word = 16'h3ccf;
			12'h3ce: tri_word = 16'h3cdf;
			12'h3cf: tri_word = 16'h3cef;
			12'h3d0: tri_word = 16'h3cff;
			12'h3d1: tri_word = 16'h3d0f;
			12'h3d2: tri_word = 16'h3d1f;
			12'h3d3: tri_word = 16'h3d2f;
			12'h3d4: tri_word = 16'h3d3f;
			12'h3d5: tri_word = 16'h3d4f;
			12'h3d6: tri_word = 16'h3d5f;
			12'h3d7: tri_word = 16'h3d6f;
			12'h3d8: tri_word = 16'h3d7f;
			12'h3d9: tri_word = 16'h3d8f;
			12'h3da: tri_word = 16'h3d9f;
			12'h3db: tri_word = 16'h3daf;
			12'h3dc: tri_word = 16'h3dbf;
			12'h3dd: tri_word = 16'h3dcf;
			12'h3de: tri_word = 16'h3ddf;
			12'h3df: tri_word = 16'h3def;
			12'h3e0: tri_word = 16'h3dff;
			12'h3e1: tri_word = 16'h3e0f;
			12'h3e2: tri_word = 16'h3e1f;
			12'h3e3: tri_word = 16'h3e2f;
			12'h3e4: tri_word = 16'h3e3f;
			12'h3e5: tri_word = 16'h3e4f;
			12'h3e6: tri_word = 16'h3e5f;
			12'h3e7: tri_word = 16'h3e6f;
			12'h3e8: tri_word = 16'h3e7f;
			12'h3e9: tri_word = 16'h3e8f;
			12'h3ea: tri_word = 16'h3e9f;
			12'h3eb: tri_word = 16'h3eaf;
			12'h3ec: tri_word = 16'h3ebf;
			12'h3ed: tri_word = 16'h3ecf;
			12'h3ee: tri_word = 16'h3edf;
			12'h3ef: tri_word = 16'h3eef;
			12'h3f0: tri_word = 16'h3eff;
			12'h3f1: tri_word = 16'h3f0f;
			12'h3f2: tri_word = 16'h3f1f;
			12'h3f3: tri_word = 16'h3f2f;
			12'h3f4: tri_word = 16'h3f3f;
			12'h3f5: tri_word = 16'h3f4f;
			12'h3f6: tri_word = 16'h3f5f;
			12'h3f7: tri_word = 16'h3f6f;
			12'h3f8: tri_word = 16'h3f7f;
			12'h3f9: tri_word = 16'h3f8f;
			12'h3fa: tri_word = 16'h3f9f;
			12'h3fb: tri_word = 16'h3faf;
			12'h3fc: tri_word = 16'h3fbf;
			12'h3fd: tri_word = 16'h3fcf;
			12'h3fe: tri_word = 16'h3fdf;
			12'h3ff: tri_word = 16'h3fef;
			12'h400: tri_word = 16'h3fff;
			12'h401: tri_word = 16'h400f;
			12'h402: tri_word = 16'h401f;
			12'h403: tri_word = 16'h402f;
			12'h404: tri_word = 16'h403f;
			12'h405: tri_word = 16'h404f;
			12'h406: tri_word = 16'h405f;
			12'h407: tri_word = 16'h406f;
			12'h408: tri_word = 16'h407f;
			12'h409: tri_word = 16'h408f;
			12'h40a: tri_word = 16'h409f;
			12'h40b: tri_word = 16'h40af;
			12'h40c: tri_word = 16'h40bf;
			12'h40d: tri_word = 16'h40cf;
			12'h40e: tri_word = 16'h40df;
			12'h40f: tri_word = 16'h40ef;
			12'h410: tri_word = 16'h40ff;
			12'h411: tri_word = 16'h410f;
			12'h412: tri_word = 16'h411f;
			12'h413: tri_word = 16'h412f;
			12'h414: tri_word = 16'h413f;
			12'h415: tri_word = 16'h414f;
			12'h416: tri_word = 16'h415f;
			12'h417: tri_word = 16'h416f;
			12'h418: tri_word = 16'h417f;
			12'h419: tri_word = 16'h418f;
			12'h41a: tri_word = 16'h419f;
			12'h41b: tri_word = 16'h41af;
			12'h41c: tri_word = 16'h41bf;
			12'h41d: tri_word = 16'h41cf;
			12'h41e: tri_word = 16'h41df;
			12'h41f: tri_word = 16'h41ef;
			12'h420: tri_word = 16'h41ff;
			12'h421: tri_word = 16'h420f;
			12'h422: tri_word = 16'h421f;
			12'h423: tri_word = 16'h422f;
			12'h424: tri_word = 16'h423f;
			12'h425: tri_word = 16'h424f;
			12'h426: tri_word = 16'h425f;
			12'h427: tri_word = 16'h426f;
			12'h428: tri_word = 16'h427f;
			12'h429: tri_word = 16'h428f;
			12'h42a: tri_word = 16'h429f;
			12'h42b: tri_word = 16'h42af;
			12'h42c: tri_word = 16'h42bf;
			12'h42d: tri_word = 16'h42cf;
			12'h42e: tri_word = 16'h42df;
			12'h42f: tri_word = 16'h42ef;
			12'h430: tri_word = 16'h42ff;
			12'h431: tri_word = 16'h430f;
			12'h432: tri_word = 16'h431f;
			12'h433: tri_word = 16'h432f;
			12'h434: tri_word = 16'h433f;
			12'h435: tri_word = 16'h434f;
			12'h436: tri_word = 16'h435f;
			12'h437: tri_word = 16'h436f;
			12'h438: tri_word = 16'h437f;
			12'h439: tri_word = 16'h438f;
			12'h43a: tri_word = 16'h439f;
			12'h43b: tri_word = 16'h43af;
			12'h43c: tri_word = 16'h43bf;
			12'h43d: tri_word = 16'h43cf;
			12'h43e: tri_word = 16'h43df;
			12'h43f: tri_word = 16'h43ef;
			12'h440: tri_word = 16'h43ff;
			12'h441: tri_word = 16'h440f;
			12'h442: tri_word = 16'h441f;
			12'h443: tri_word = 16'h442f;
			12'h444: tri_word = 16'h443f;
			12'h445: tri_word = 16'h444f;
			12'h446: tri_word = 16'h445f;
			12'h447: tri_word = 16'h446f;
			12'h448: tri_word = 16'h447f;
			12'h449: tri_word = 16'h448f;
			12'h44a: tri_word = 16'h449f;
			12'h44b: tri_word = 16'h44af;
			12'h44c: tri_word = 16'h44bf;
			12'h44d: tri_word = 16'h44cf;
			12'h44e: tri_word = 16'h44df;
			12'h44f: tri_word = 16'h44ef;
			12'h450: tri_word = 16'h44ff;
			12'h451: tri_word = 16'h450f;
			12'h452: tri_word = 16'h451f;
			12'h453: tri_word = 16'h452f;
			12'h454: tri_word = 16'h453f;
			12'h455: tri_word = 16'h454f;
			12'h456: tri_word = 16'h455f;
			12'h457: tri_word = 16'h456f;
			12'h458: tri_word = 16'h457f;
			12'h459: tri_word = 16'h458f;
			12'h45a: tri_word = 16'h459f;
			12'h45b: tri_word = 16'h45af;
			12'h45c: tri_word = 16'h45bf;
			12'h45d: tri_word = 16'h45cf;
			12'h45e: tri_word = 16'h45df;
			12'h45f: tri_word = 16'h45ef;
			12'h460: tri_word = 16'h45ff;
			12'h461: tri_word = 16'h460f;
			12'h462: tri_word = 16'h461f;
			12'h463: tri_word = 16'h462f;
			12'h464: tri_word = 16'h463f;
			12'h465: tri_word = 16'h464f;
			12'h466: tri_word = 16'h465f;
			12'h467: tri_word = 16'h466f;
			12'h468: tri_word = 16'h467f;
			12'h469: tri_word = 16'h468f;
			12'h46a: tri_word = 16'h469f;
			12'h46b: tri_word = 16'h46af;
			12'h46c: tri_word = 16'h46bf;
			12'h46d: tri_word = 16'h46cf;
			12'h46e: tri_word = 16'h46df;
			12'h46f: tri_word = 16'h46ef;
			12'h470: tri_word = 16'h46ff;
			12'h471: tri_word = 16'h470f;
			12'h472: tri_word = 16'h471f;
			12'h473: tri_word = 16'h472f;
			12'h474: tri_word = 16'h473f;
			12'h475: tri_word = 16'h474f;
			12'h476: tri_word = 16'h475f;
			12'h477: tri_word = 16'h476f;
			12'h478: tri_word = 16'h477f;
			12'h479: tri_word = 16'h478f;
			12'h47a: tri_word = 16'h479f;
			12'h47b: tri_word = 16'h47af;
			12'h47c: tri_word = 16'h47bf;
			12'h47d: tri_word = 16'h47cf;
			12'h47e: tri_word = 16'h47df;
			12'h47f: tri_word = 16'h47ef;
			12'h480: tri_word = 16'h47ff;
			12'h481: tri_word = 16'h480f;
			12'h482: tri_word = 16'h481f;
			12'h483: tri_word = 16'h482f;
			12'h484: tri_word = 16'h483f;
			12'h485: tri_word = 16'h484f;
			12'h486: tri_word = 16'h485f;
			12'h487: tri_word = 16'h486f;
			12'h488: tri_word = 16'h487f;
			12'h489: tri_word = 16'h488f;
			12'h48a: tri_word = 16'h489f;
			12'h48b: tri_word = 16'h48af;
			12'h48c: tri_word = 16'h48bf;
			12'h48d: tri_word = 16'h48cf;
			12'h48e: tri_word = 16'h48df;
			12'h48f: tri_word = 16'h48ef;
			12'h490: tri_word = 16'h48ff;
			12'h491: tri_word = 16'h490f;
			12'h492: tri_word = 16'h491f;
			12'h493: tri_word = 16'h492f;
			12'h494: tri_word = 16'h493f;
			12'h495: tri_word = 16'h494f;
			12'h496: tri_word = 16'h495f;
			12'h497: tri_word = 16'h496f;
			12'h498: tri_word = 16'h497f;
			12'h499: tri_word = 16'h498f;
			12'h49a: tri_word = 16'h499f;
			12'h49b: tri_word = 16'h49af;
			12'h49c: tri_word = 16'h49bf;
			12'h49d: tri_word = 16'h49cf;
			12'h49e: tri_word = 16'h49df;
			12'h49f: tri_word = 16'h49ef;
			12'h4a0: tri_word = 16'h49ff;
			12'h4a1: tri_word = 16'h4a0f;
			12'h4a2: tri_word = 16'h4a1f;
			12'h4a3: tri_word = 16'h4a2f;
			12'h4a4: tri_word = 16'h4a3f;
			12'h4a5: tri_word = 16'h4a4f;
			12'h4a6: tri_word = 16'h4a5f;
			12'h4a7: tri_word = 16'h4a6f;
			12'h4a8: tri_word = 16'h4a7f;
			12'h4a9: tri_word = 16'h4a8f;
			12'h4aa: tri_word = 16'h4a9f;
			12'h4ab: tri_word = 16'h4aaf;
			12'h4ac: tri_word = 16'h4abf;
			12'h4ad: tri_word = 16'h4acf;
			12'h4ae: tri_word = 16'h4adf;
			12'h4af: tri_word = 16'h4aef;
			12'h4b0: tri_word = 16'h4aff;
			12'h4b1: tri_word = 16'h4b0f;
			12'h4b2: tri_word = 16'h4b1f;
			12'h4b3: tri_word = 16'h4b2f;
			12'h4b4: tri_word = 16'h4b3f;
			12'h4b5: tri_word = 16'h4b4f;
			12'h4b6: tri_word = 16'h4b5f;
			12'h4b7: tri_word = 16'h4b6f;
			12'h4b8: tri_word = 16'h4b7f;
			12'h4b9: tri_word = 16'h4b8f;
			12'h4ba: tri_word = 16'h4b9f;
			12'h4bb: tri_word = 16'h4baf;
			12'h4bc: tri_word = 16'h4bbf;
			12'h4bd: tri_word = 16'h4bcf;
			12'h4be: tri_word = 16'h4bdf;
			12'h4bf: tri_word = 16'h4bef;
			12'h4c0: tri_word = 16'h4bff;
			12'h4c1: tri_word = 16'h4c0f;
			12'h4c2: tri_word = 16'h4c1f;
			12'h4c3: tri_word = 16'h4c2f;
			12'h4c4: tri_word = 16'h4c3f;
			12'h4c5: tri_word = 16'h4c4f;
			12'h4c6: tri_word = 16'h4c5f;
			12'h4c7: tri_word = 16'h4c6f;
			12'h4c8: tri_word = 16'h4c7f;
			12'h4c9: tri_word = 16'h4c8f;
			12'h4ca: tri_word = 16'h4c9f;
			12'h4cb: tri_word = 16'h4caf;
			12'h4cc: tri_word = 16'h4cbf;
			12'h4cd: tri_word = 16'h4ccf;
			12'h4ce: tri_word = 16'h4cdf;
			12'h4cf: tri_word = 16'h4cef;
			12'h4d0: tri_word = 16'h4cff;
			12'h4d1: tri_word = 16'h4d0f;
			12'h4d2: tri_word = 16'h4d1f;
			12'h4d3: tri_word = 16'h4d2f;
			12'h4d4: tri_word = 16'h4d3f;
			12'h4d5: tri_word = 16'h4d4f;
			12'h4d6: tri_word = 16'h4d5f;
			12'h4d7: tri_word = 16'h4d6f;
			12'h4d8: tri_word = 16'h4d7f;
			12'h4d9: tri_word = 16'h4d8f;
			12'h4da: tri_word = 16'h4d9f;
			12'h4db: tri_word = 16'h4daf;
			12'h4dc: tri_word = 16'h4dbf;
			12'h4dd: tri_word = 16'h4dcf;
			12'h4de: tri_word = 16'h4ddf;
			12'h4df: tri_word = 16'h4def;
			12'h4e0: tri_word = 16'h4dff;
			12'h4e1: tri_word = 16'h4e0f;
			12'h4e2: tri_word = 16'h4e1f;
			12'h4e3: tri_word = 16'h4e2f;
			12'h4e4: tri_word = 16'h4e3f;
			12'h4e5: tri_word = 16'h4e4f;
			12'h4e6: tri_word = 16'h4e5f;
			12'h4e7: tri_word = 16'h4e6f;
			12'h4e8: tri_word = 16'h4e7f;
			12'h4e9: tri_word = 16'h4e8f;
			12'h4ea: tri_word = 16'h4e9f;
			12'h4eb: tri_word = 16'h4eaf;
			12'h4ec: tri_word = 16'h4ebf;
			12'h4ed: tri_word = 16'h4ecf;
			12'h4ee: tri_word = 16'h4edf;
			12'h4ef: tri_word = 16'h4eef;
			12'h4f0: tri_word = 16'h4eff;
			12'h4f1: tri_word = 16'h4f0f;
			12'h4f2: tri_word = 16'h4f1f;
			12'h4f3: tri_word = 16'h4f2f;
			12'h4f4: tri_word = 16'h4f3f;
			12'h4f5: tri_word = 16'h4f4f;
			12'h4f6: tri_word = 16'h4f5f;
			12'h4f7: tri_word = 16'h4f6f;
			12'h4f8: tri_word = 16'h4f7f;
			12'h4f9: tri_word = 16'h4f8f;
			12'h4fa: tri_word = 16'h4f9f;
			12'h4fb: tri_word = 16'h4faf;
			12'h4fc: tri_word = 16'h4fbf;
			12'h4fd: tri_word = 16'h4fcf;
			12'h4fe: tri_word = 16'h4fdf;
			12'h4ff: tri_word = 16'h4fef;
			12'h500: tri_word = 16'h4fff;
			12'h501: tri_word = 16'h500f;
			12'h502: tri_word = 16'h501f;
			12'h503: tri_word = 16'h502f;
			12'h504: tri_word = 16'h503f;
			12'h505: tri_word = 16'h504f;
			12'h506: tri_word = 16'h505f;
			12'h507: tri_word = 16'h506f;
			12'h508: tri_word = 16'h507f;
			12'h509: tri_word = 16'h508f;
			12'h50a: tri_word = 16'h509f;
			12'h50b: tri_word = 16'h50af;
			12'h50c: tri_word = 16'h50bf;
			12'h50d: tri_word = 16'h50cf;
			12'h50e: tri_word = 16'h50df;
			12'h50f: tri_word = 16'h50ef;
			12'h510: tri_word = 16'h50ff;
			12'h511: tri_word = 16'h510f;
			12'h512: tri_word = 16'h511f;
			12'h513: tri_word = 16'h512f;
			12'h514: tri_word = 16'h513f;
			12'h515: tri_word = 16'h514f;
			12'h516: tri_word = 16'h515f;
			12'h517: tri_word = 16'h516f;
			12'h518: tri_word = 16'h517f;
			12'h519: tri_word = 16'h518f;
			12'h51a: tri_word = 16'h519f;
			12'h51b: tri_word = 16'h51af;
			12'h51c: tri_word = 16'h51bf;
			12'h51d: tri_word = 16'h51cf;
			12'h51e: tri_word = 16'h51df;
			12'h51f: tri_word = 16'h51ef;
			12'h520: tri_word = 16'h51ff;
			12'h521: tri_word = 16'h520f;
			12'h522: tri_word = 16'h521f;
			12'h523: tri_word = 16'h522f;
			12'h524: tri_word = 16'h523f;
			12'h525: tri_word = 16'h524f;
			12'h526: tri_word = 16'h525f;
			12'h527: tri_word = 16'h526f;
			12'h528: tri_word = 16'h527f;
			12'h529: tri_word = 16'h528f;
			12'h52a: tri_word = 16'h529f;
			12'h52b: tri_word = 16'h52af;
			12'h52c: tri_word = 16'h52bf;
			12'h52d: tri_word = 16'h52cf;
			12'h52e: tri_word = 16'h52df;
			12'h52f: tri_word = 16'h52ef;
			12'h530: tri_word = 16'h52ff;
			12'h531: tri_word = 16'h530f;
			12'h532: tri_word = 16'h531f;
			12'h533: tri_word = 16'h532f;
			12'h534: tri_word = 16'h533f;
			12'h535: tri_word = 16'h534f;
			12'h536: tri_word = 16'h535f;
			12'h537: tri_word = 16'h536f;
			12'h538: tri_word = 16'h537f;
			12'h539: tri_word = 16'h538f;
			12'h53a: tri_word = 16'h539f;
			12'h53b: tri_word = 16'h53af;
			12'h53c: tri_word = 16'h53bf;
			12'h53d: tri_word = 16'h53cf;
			12'h53e: tri_word = 16'h53df;
			12'h53f: tri_word = 16'h53ef;
			12'h540: tri_word = 16'h53ff;
			12'h541: tri_word = 16'h540f;
			12'h542: tri_word = 16'h541f;
			12'h543: tri_word = 16'h542f;
			12'h544: tri_word = 16'h543f;
			12'h545: tri_word = 16'h544f;
			12'h546: tri_word = 16'h545f;
			12'h547: tri_word = 16'h546f;
			12'h548: tri_word = 16'h547f;
			12'h549: tri_word = 16'h548f;
			12'h54a: tri_word = 16'h549f;
			12'h54b: tri_word = 16'h54af;
			12'h54c: tri_word = 16'h54bf;
			12'h54d: tri_word = 16'h54cf;
			12'h54e: tri_word = 16'h54df;
			12'h54f: tri_word = 16'h54ef;
			12'h550: tri_word = 16'h54ff;
			12'h551: tri_word = 16'h550f;
			12'h552: tri_word = 16'h551f;
			12'h553: tri_word = 16'h552f;
			12'h554: tri_word = 16'h553f;
			12'h555: tri_word = 16'h554f;
			12'h556: tri_word = 16'h555f;
			12'h557: tri_word = 16'h556f;
			12'h558: tri_word = 16'h557f;
			12'h559: tri_word = 16'h558f;
			12'h55a: tri_word = 16'h559f;
			12'h55b: tri_word = 16'h55af;
			12'h55c: tri_word = 16'h55bf;
			12'h55d: tri_word = 16'h55cf;
			12'h55e: tri_word = 16'h55df;
			12'h55f: tri_word = 16'h55ef;
			12'h560: tri_word = 16'h55ff;
			12'h561: tri_word = 16'h560f;
			12'h562: tri_word = 16'h561f;
			12'h563: tri_word = 16'h562f;
			12'h564: tri_word = 16'h563f;
			12'h565: tri_word = 16'h564f;
			12'h566: tri_word = 16'h565f;
			12'h567: tri_word = 16'h566f;
			12'h568: tri_word = 16'h567f;
			12'h569: tri_word = 16'h568f;
			12'h56a: tri_word = 16'h569f;
			12'h56b: tri_word = 16'h56af;
			12'h56c: tri_word = 16'h56bf;
			12'h56d: tri_word = 16'h56cf;
			12'h56e: tri_word = 16'h56df;
			12'h56f: tri_word = 16'h56ef;
			12'h570: tri_word = 16'h56ff;
			12'h571: tri_word = 16'h570f;
			12'h572: tri_word = 16'h571f;
			12'h573: tri_word = 16'h572f;
			12'h574: tri_word = 16'h573f;
			12'h575: tri_word = 16'h574f;
			12'h576: tri_word = 16'h575f;
			12'h577: tri_word = 16'h576f;
			12'h578: tri_word = 16'h577f;
			12'h579: tri_word = 16'h578f;
			12'h57a: tri_word = 16'h579f;
			12'h57b: tri_word = 16'h57af;
			12'h57c: tri_word = 16'h57bf;
			12'h57d: tri_word = 16'h57cf;
			12'h57e: tri_word = 16'h57df;
			12'h57f: tri_word = 16'h57ef;
			12'h580: tri_word = 16'h57ff;
			12'h581: tri_word = 16'h580f;
			12'h582: tri_word = 16'h581f;
			12'h583: tri_word = 16'h582f;
			12'h584: tri_word = 16'h583f;
			12'h585: tri_word = 16'h584f;
			12'h586: tri_word = 16'h585f;
			12'h587: tri_word = 16'h586f;
			12'h588: tri_word = 16'h587f;
			12'h589: tri_word = 16'h588f;
			12'h58a: tri_word = 16'h589f;
			12'h58b: tri_word = 16'h58af;
			12'h58c: tri_word = 16'h58bf;
			12'h58d: tri_word = 16'h58cf;
			12'h58e: tri_word = 16'h58df;
			12'h58f: tri_word = 16'h58ef;
			12'h590: tri_word = 16'h58ff;
			12'h591: tri_word = 16'h590f;
			12'h592: tri_word = 16'h591f;
			12'h593: tri_word = 16'h592f;
			12'h594: tri_word = 16'h593f;
			12'h595: tri_word = 16'h594f;
			12'h596: tri_word = 16'h595f;
			12'h597: tri_word = 16'h596f;
			12'h598: tri_word = 16'h597f;
			12'h599: tri_word = 16'h598f;
			12'h59a: tri_word = 16'h599f;
			12'h59b: tri_word = 16'h59af;
			12'h59c: tri_word = 16'h59bf;
			12'h59d: tri_word = 16'h59cf;
			12'h59e: tri_word = 16'h59df;
			12'h59f: tri_word = 16'h59ef;
			12'h5a0: tri_word = 16'h59ff;
			12'h5a1: tri_word = 16'h5a0f;
			12'h5a2: tri_word = 16'h5a1f;
			12'h5a3: tri_word = 16'h5a2f;
			12'h5a4: tri_word = 16'h5a3f;
			12'h5a5: tri_word = 16'h5a4f;
			12'h5a6: tri_word = 16'h5a5f;
			12'h5a7: tri_word = 16'h5a6f;
			12'h5a8: tri_word = 16'h5a7f;
			12'h5a9: tri_word = 16'h5a8f;
			12'h5aa: tri_word = 16'h5a9f;
			12'h5ab: tri_word = 16'h5aaf;
			12'h5ac: tri_word = 16'h5abf;
			12'h5ad: tri_word = 16'h5acf;
			12'h5ae: tri_word = 16'h5adf;
			12'h5af: tri_word = 16'h5aef;
			12'h5b0: tri_word = 16'h5aff;
			12'h5b1: tri_word = 16'h5b0f;
			12'h5b2: tri_word = 16'h5b1f;
			12'h5b3: tri_word = 16'h5b2f;
			12'h5b4: tri_word = 16'h5b3f;
			12'h5b5: tri_word = 16'h5b4f;
			12'h5b6: tri_word = 16'h5b5f;
			12'h5b7: tri_word = 16'h5b6f;
			12'h5b8: tri_word = 16'h5b7f;
			12'h5b9: tri_word = 16'h5b8f;
			12'h5ba: tri_word = 16'h5b9f;
			12'h5bb: tri_word = 16'h5baf;
			12'h5bc: tri_word = 16'h5bbf;
			12'h5bd: tri_word = 16'h5bcf;
			12'h5be: tri_word = 16'h5bdf;
			12'h5bf: tri_word = 16'h5bef;
			12'h5c0: tri_word = 16'h5bff;
			12'h5c1: tri_word = 16'h5c0f;
			12'h5c2: tri_word = 16'h5c1f;
			12'h5c3: tri_word = 16'h5c2f;
			12'h5c4: tri_word = 16'h5c3f;
			12'h5c5: tri_word = 16'h5c4f;
			12'h5c6: tri_word = 16'h5c5f;
			12'h5c7: tri_word = 16'h5c6f;
			12'h5c8: tri_word = 16'h5c7f;
			12'h5c9: tri_word = 16'h5c8f;
			12'h5ca: tri_word = 16'h5c9f;
			12'h5cb: tri_word = 16'h5caf;
			12'h5cc: tri_word = 16'h5cbf;
			12'h5cd: tri_word = 16'h5ccf;
			12'h5ce: tri_word = 16'h5cdf;
			12'h5cf: tri_word = 16'h5cef;
			12'h5d0: tri_word = 16'h5cff;
			12'h5d1: tri_word = 16'h5d0f;
			12'h5d2: tri_word = 16'h5d1f;
			12'h5d3: tri_word = 16'h5d2f;
			12'h5d4: tri_word = 16'h5d3f;
			12'h5d5: tri_word = 16'h5d4f;
			12'h5d6: tri_word = 16'h5d5f;
			12'h5d7: tri_word = 16'h5d6f;
			12'h5d8: tri_word = 16'h5d7f;
			12'h5d9: tri_word = 16'h5d8f;
			12'h5da: tri_word = 16'h5d9f;
			12'h5db: tri_word = 16'h5daf;
			12'h5dc: tri_word = 16'h5dbf;
			12'h5dd: tri_word = 16'h5dcf;
			12'h5de: tri_word = 16'h5ddf;
			12'h5df: tri_word = 16'h5def;
			12'h5e0: tri_word = 16'h5dff;
			12'h5e1: tri_word = 16'h5e0f;
			12'h5e2: tri_word = 16'h5e1f;
			12'h5e3: tri_word = 16'h5e2f;
			12'h5e4: tri_word = 16'h5e3f;
			12'h5e5: tri_word = 16'h5e4f;
			12'h5e6: tri_word = 16'h5e5f;
			12'h5e7: tri_word = 16'h5e6f;
			12'h5e8: tri_word = 16'h5e7f;
			12'h5e9: tri_word = 16'h5e8f;
			12'h5ea: tri_word = 16'h5e9f;
			12'h5eb: tri_word = 16'h5eaf;
			12'h5ec: tri_word = 16'h5ebf;
			12'h5ed: tri_word = 16'h5ecf;
			12'h5ee: tri_word = 16'h5edf;
			12'h5ef: tri_word = 16'h5eef;
			12'h5f0: tri_word = 16'h5eff;
			12'h5f1: tri_word = 16'h5f0f;
			12'h5f2: tri_word = 16'h5f1f;
			12'h5f3: tri_word = 16'h5f2f;
			12'h5f4: tri_word = 16'h5f3f;
			12'h5f5: tri_word = 16'h5f4f;
			12'h5f6: tri_word = 16'h5f5f;
			12'h5f7: tri_word = 16'h5f6f;
			12'h5f8: tri_word = 16'h5f7f;
			12'h5f9: tri_word = 16'h5f8f;
			12'h5fa: tri_word = 16'h5f9f;
			12'h5fb: tri_word = 16'h5faf;
			12'h5fc: tri_word = 16'h5fbf;
			12'h5fd: tri_word = 16'h5fcf;
			12'h5fe: tri_word = 16'h5fdf;
			12'h5ff: tri_word = 16'h5fef;
			12'h600: tri_word = 16'h5fff;
			12'h601: tri_word = 16'h600f;
			12'h602: tri_word = 16'h601f;
			12'h603: tri_word = 16'h602f;
			12'h604: tri_word = 16'h603f;
			12'h605: tri_word = 16'h604f;
			12'h606: tri_word = 16'h605f;
			12'h607: tri_word = 16'h606f;
			12'h608: tri_word = 16'h607f;
			12'h609: tri_word = 16'h608f;
			12'h60a: tri_word = 16'h609f;
			12'h60b: tri_word = 16'h60af;
			12'h60c: tri_word = 16'h60bf;
			12'h60d: tri_word = 16'h60cf;
			12'h60e: tri_word = 16'h60df;
			12'h60f: tri_word = 16'h60ef;
			12'h610: tri_word = 16'h60ff;
			12'h611: tri_word = 16'h610f;
			12'h612: tri_word = 16'h611f;
			12'h613: tri_word = 16'h612f;
			12'h614: tri_word = 16'h613f;
			12'h615: tri_word = 16'h614f;
			12'h616: tri_word = 16'h615f;
			12'h617: tri_word = 16'h616f;
			12'h618: tri_word = 16'h617f;
			12'h619: tri_word = 16'h618f;
			12'h61a: tri_word = 16'h619f;
			12'h61b: tri_word = 16'h61af;
			12'h61c: tri_word = 16'h61bf;
			12'h61d: tri_word = 16'h61cf;
			12'h61e: tri_word = 16'h61df;
			12'h61f: tri_word = 16'h61ef;
			12'h620: tri_word = 16'h61ff;
			12'h621: tri_word = 16'h620f;
			12'h622: tri_word = 16'h621f;
			12'h623: tri_word = 16'h622f;
			12'h624: tri_word = 16'h623f;
			12'h625: tri_word = 16'h624f;
			12'h626: tri_word = 16'h625f;
			12'h627: tri_word = 16'h626f;
			12'h628: tri_word = 16'h627f;
			12'h629: tri_word = 16'h628f;
			12'h62a: tri_word = 16'h629f;
			12'h62b: tri_word = 16'h62af;
			12'h62c: tri_word = 16'h62bf;
			12'h62d: tri_word = 16'h62cf;
			12'h62e: tri_word = 16'h62df;
			12'h62f: tri_word = 16'h62ef;
			12'h630: tri_word = 16'h62ff;
			12'h631: tri_word = 16'h630f;
			12'h632: tri_word = 16'h631f;
			12'h633: tri_word = 16'h632f;
			12'h634: tri_word = 16'h633f;
			12'h635: tri_word = 16'h634f;
			12'h636: tri_word = 16'h635f;
			12'h637: tri_word = 16'h636f;
			12'h638: tri_word = 16'h637f;
			12'h639: tri_word = 16'h638f;
			12'h63a: tri_word = 16'h639f;
			12'h63b: tri_word = 16'h63af;
			12'h63c: tri_word = 16'h63bf;
			12'h63d: tri_word = 16'h63cf;
			12'h63e: tri_word = 16'h63df;
			12'h63f: tri_word = 16'h63ef;
			12'h640: tri_word = 16'h63ff;
			12'h641: tri_word = 16'h640f;
			12'h642: tri_word = 16'h641f;
			12'h643: tri_word = 16'h642f;
			12'h644: tri_word = 16'h643f;
			12'h645: tri_word = 16'h644f;
			12'h646: tri_word = 16'h645f;
			12'h647: tri_word = 16'h646f;
			12'h648: tri_word = 16'h647f;
			12'h649: tri_word = 16'h648f;
			12'h64a: tri_word = 16'h649f;
			12'h64b: tri_word = 16'h64af;
			12'h64c: tri_word = 16'h64bf;
			12'h64d: tri_word = 16'h64cf;
			12'h64e: tri_word = 16'h64df;
			12'h64f: tri_word = 16'h64ef;
			12'h650: tri_word = 16'h64ff;
			12'h651: tri_word = 16'h650f;
			12'h652: tri_word = 16'h651f;
			12'h653: tri_word = 16'h652f;
			12'h654: tri_word = 16'h653f;
			12'h655: tri_word = 16'h654f;
			12'h656: tri_word = 16'h655f;
			12'h657: tri_word = 16'h656f;
			12'h658: tri_word = 16'h657f;
			12'h659: tri_word = 16'h658f;
			12'h65a: tri_word = 16'h659f;
			12'h65b: tri_word = 16'h65af;
			12'h65c: tri_word = 16'h65bf;
			12'h65d: tri_word = 16'h65cf;
			12'h65e: tri_word = 16'h65df;
			12'h65f: tri_word = 16'h65ef;
			12'h660: tri_word = 16'h65ff;
			12'h661: tri_word = 16'h660f;
			12'h662: tri_word = 16'h661f;
			12'h663: tri_word = 16'h662f;
			12'h664: tri_word = 16'h663f;
			12'h665: tri_word = 16'h664f;
			12'h666: tri_word = 16'h665f;
			12'h667: tri_word = 16'h666f;
			12'h668: tri_word = 16'h667f;
			12'h669: tri_word = 16'h668f;
			12'h66a: tri_word = 16'h669f;
			12'h66b: tri_word = 16'h66af;
			12'h66c: tri_word = 16'h66bf;
			12'h66d: tri_word = 16'h66cf;
			12'h66e: tri_word = 16'h66df;
			12'h66f: tri_word = 16'h66ef;
			12'h670: tri_word = 16'h66ff;
			12'h671: tri_word = 16'h670f;
			12'h672: tri_word = 16'h671f;
			12'h673: tri_word = 16'h672f;
			12'h674: tri_word = 16'h673f;
			12'h675: tri_word = 16'h674f;
			12'h676: tri_word = 16'h675f;
			12'h677: tri_word = 16'h676f;
			12'h678: tri_word = 16'h677f;
			12'h679: tri_word = 16'h678f;
			12'h67a: tri_word = 16'h679f;
			12'h67b: tri_word = 16'h67af;
			12'h67c: tri_word = 16'h67bf;
			12'h67d: tri_word = 16'h67cf;
			12'h67e: tri_word = 16'h67df;
			12'h67f: tri_word = 16'h67ef;
			12'h680: tri_word = 16'h67ff;
			12'h681: tri_word = 16'h680f;
			12'h682: tri_word = 16'h681f;
			12'h683: tri_word = 16'h682f;
			12'h684: tri_word = 16'h683f;
			12'h685: tri_word = 16'h684f;
			12'h686: tri_word = 16'h685f;
			12'h687: tri_word = 16'h686f;
			12'h688: tri_word = 16'h687f;
			12'h689: tri_word = 16'h688f;
			12'h68a: tri_word = 16'h689f;
			12'h68b: tri_word = 16'h68af;
			12'h68c: tri_word = 16'h68bf;
			12'h68d: tri_word = 16'h68cf;
			12'h68e: tri_word = 16'h68df;
			12'h68f: tri_word = 16'h68ef;
			12'h690: tri_word = 16'h68ff;
			12'h691: tri_word = 16'h690f;
			12'h692: tri_word = 16'h691f;
			12'h693: tri_word = 16'h692f;
			12'h694: tri_word = 16'h693f;
			12'h695: tri_word = 16'h694f;
			12'h696: tri_word = 16'h695f;
			12'h697: tri_word = 16'h696f;
			12'h698: tri_word = 16'h697f;
			12'h699: tri_word = 16'h698f;
			12'h69a: tri_word = 16'h699f;
			12'h69b: tri_word = 16'h69af;
			12'h69c: tri_word = 16'h69bf;
			12'h69d: tri_word = 16'h69cf;
			12'h69e: tri_word = 16'h69df;
			12'h69f: tri_word = 16'h69ef;
			12'h6a0: tri_word = 16'h69ff;
			12'h6a1: tri_word = 16'h6a0f;
			12'h6a2: tri_word = 16'h6a1f;
			12'h6a3: tri_word = 16'h6a2f;
			12'h6a4: tri_word = 16'h6a3f;
			12'h6a5: tri_word = 16'h6a4f;
			12'h6a6: tri_word = 16'h6a5f;
			12'h6a7: tri_word = 16'h6a6f;
			12'h6a8: tri_word = 16'h6a7f;
			12'h6a9: tri_word = 16'h6a8f;
			12'h6aa: tri_word = 16'h6a9f;
			12'h6ab: tri_word = 16'h6aaf;
			12'h6ac: tri_word = 16'h6abf;
			12'h6ad: tri_word = 16'h6acf;
			12'h6ae: tri_word = 16'h6adf;
			12'h6af: tri_word = 16'h6aef;
			12'h6b0: tri_word = 16'h6aff;
			12'h6b1: tri_word = 16'h6b0f;
			12'h6b2: tri_word = 16'h6b1f;
			12'h6b3: tri_word = 16'h6b2f;
			12'h6b4: tri_word = 16'h6b3f;
			12'h6b5: tri_word = 16'h6b4f;
			12'h6b6: tri_word = 16'h6b5f;
			12'h6b7: tri_word = 16'h6b6f;
			12'h6b8: tri_word = 16'h6b7f;
			12'h6b9: tri_word = 16'h6b8f;
			12'h6ba: tri_word = 16'h6b9f;
			12'h6bb: tri_word = 16'h6baf;
			12'h6bc: tri_word = 16'h6bbf;
			12'h6bd: tri_word = 16'h6bcf;
			12'h6be: tri_word = 16'h6bdf;
			12'h6bf: tri_word = 16'h6bef;
			12'h6c0: tri_word = 16'h6bff;
			12'h6c1: tri_word = 16'h6c0f;
			12'h6c2: tri_word = 16'h6c1f;
			12'h6c3: tri_word = 16'h6c2f;
			12'h6c4: tri_word = 16'h6c3f;
			12'h6c5: tri_word = 16'h6c4f;
			12'h6c6: tri_word = 16'h6c5f;
			12'h6c7: tri_word = 16'h6c6f;
			12'h6c8: tri_word = 16'h6c7f;
			12'h6c9: tri_word = 16'h6c8f;
			12'h6ca: tri_word = 16'h6c9f;
			12'h6cb: tri_word = 16'h6caf;
			12'h6cc: tri_word = 16'h6cbf;
			12'h6cd: tri_word = 16'h6ccf;
			12'h6ce: tri_word = 16'h6cdf;
			12'h6cf: tri_word = 16'h6cef;
			12'h6d0: tri_word = 16'h6cff;
			12'h6d1: tri_word = 16'h6d0f;
			12'h6d2: tri_word = 16'h6d1f;
			12'h6d3: tri_word = 16'h6d2f;
			12'h6d4: tri_word = 16'h6d3f;
			12'h6d5: tri_word = 16'h6d4f;
			12'h6d6: tri_word = 16'h6d5f;
			12'h6d7: tri_word = 16'h6d6f;
			12'h6d8: tri_word = 16'h6d7f;
			12'h6d9: tri_word = 16'h6d8f;
			12'h6da: tri_word = 16'h6d9f;
			12'h6db: tri_word = 16'h6daf;
			12'h6dc: tri_word = 16'h6dbf;
			12'h6dd: tri_word = 16'h6dcf;
			12'h6de: tri_word = 16'h6ddf;
			12'h6df: tri_word = 16'h6def;
			12'h6e0: tri_word = 16'h6dff;
			12'h6e1: tri_word = 16'h6e0f;
			12'h6e2: tri_word = 16'h6e1f;
			12'h6e3: tri_word = 16'h6e2f;
			12'h6e4: tri_word = 16'h6e3f;
			12'h6e5: tri_word = 16'h6e4f;
			12'h6e6: tri_word = 16'h6e5f;
			12'h6e7: tri_word = 16'h6e6f;
			12'h6e8: tri_word = 16'h6e7f;
			12'h6e9: tri_word = 16'h6e8f;
			12'h6ea: tri_word = 16'h6e9f;
			12'h6eb: tri_word = 16'h6eaf;
			12'h6ec: tri_word = 16'h6ebf;
			12'h6ed: tri_word = 16'h6ecf;
			12'h6ee: tri_word = 16'h6edf;
			12'h6ef: tri_word = 16'h6eef;
			12'h6f0: tri_word = 16'h6eff;
			12'h6f1: tri_word = 16'h6f0f;
			12'h6f2: tri_word = 16'h6f1f;
			12'h6f3: tri_word = 16'h6f2f;
			12'h6f4: tri_word = 16'h6f3f;
			12'h6f5: tri_word = 16'h6f4f;
			12'h6f6: tri_word = 16'h6f5f;
			12'h6f7: tri_word = 16'h6f6f;
			12'h6f8: tri_word = 16'h6f7f;
			12'h6f9: tri_word = 16'h6f8f;
			12'h6fa: tri_word = 16'h6f9f;
			12'h6fb: tri_word = 16'h6faf;
			12'h6fc: tri_word = 16'h6fbf;
			12'h6fd: tri_word = 16'h6fcf;
			12'h6fe: tri_word = 16'h6fdf;
			12'h6ff: tri_word = 16'h6fef;
			12'h700: tri_word = 16'h6fff;
			12'h701: tri_word = 16'h700f;
			12'h702: tri_word = 16'h701f;
			12'h703: tri_word = 16'h702f;
			12'h704: tri_word = 16'h703f;
			12'h705: tri_word = 16'h704f;
			12'h706: tri_word = 16'h705f;
			12'h707: tri_word = 16'h706f;
			12'h708: tri_word = 16'h707f;
			12'h709: tri_word = 16'h708f;
			12'h70a: tri_word = 16'h709f;
			12'h70b: tri_word = 16'h70af;
			12'h70c: tri_word = 16'h70bf;
			12'h70d: tri_word = 16'h70cf;
			12'h70e: tri_word = 16'h70df;
			12'h70f: tri_word = 16'h70ef;
			12'h710: tri_word = 16'h70ff;
			12'h711: tri_word = 16'h710f;
			12'h712: tri_word = 16'h711f;
			12'h713: tri_word = 16'h712f;
			12'h714: tri_word = 16'h713f;
			12'h715: tri_word = 16'h714f;
			12'h716: tri_word = 16'h715f;
			12'h717: tri_word = 16'h716f;
			12'h718: tri_word = 16'h717f;
			12'h719: tri_word = 16'h718f;
			12'h71a: tri_word = 16'h719f;
			12'h71b: tri_word = 16'h71af;
			12'h71c: tri_word = 16'h71bf;
			12'h71d: tri_word = 16'h71cf;
			12'h71e: tri_word = 16'h71df;
			12'h71f: tri_word = 16'h71ef;
			12'h720: tri_word = 16'h71ff;
			12'h721: tri_word = 16'h720f;
			12'h722: tri_word = 16'h721f;
			12'h723: tri_word = 16'h722f;
			12'h724: tri_word = 16'h723f;
			12'h725: tri_word = 16'h724f;
			12'h726: tri_word = 16'h725f;
			12'h727: tri_word = 16'h726f;
			12'h728: tri_word = 16'h727f;
			12'h729: tri_word = 16'h728f;
			12'h72a: tri_word = 16'h729f;
			12'h72b: tri_word = 16'h72af;
			12'h72c: tri_word = 16'h72bf;
			12'h72d: tri_word = 16'h72cf;
			12'h72e: tri_word = 16'h72df;
			12'h72f: tri_word = 16'h72ef;
			12'h730: tri_word = 16'h72ff;
			12'h731: tri_word = 16'h730f;
			12'h732: tri_word = 16'h731f;
			12'h733: tri_word = 16'h732f;
			12'h734: tri_word = 16'h733f;
			12'h735: tri_word = 16'h734f;
			12'h736: tri_word = 16'h735f;
			12'h737: tri_word = 16'h736f;
			12'h738: tri_word = 16'h737f;
			12'h739: tri_word = 16'h738f;
			12'h73a: tri_word = 16'h739f;
			12'h73b: tri_word = 16'h73af;
			12'h73c: tri_word = 16'h73bf;
			12'h73d: tri_word = 16'h73cf;
			12'h73e: tri_word = 16'h73df;
			12'h73f: tri_word = 16'h73ef;
			12'h740: tri_word = 16'h73ff;
			12'h741: tri_word = 16'h740f;
			12'h742: tri_word = 16'h741f;
			12'h743: tri_word = 16'h742f;
			12'h744: tri_word = 16'h743f;
			12'h745: tri_word = 16'h744f;
			12'h746: tri_word = 16'h745f;
			12'h747: tri_word = 16'h746f;
			12'h748: tri_word = 16'h747f;
			12'h749: tri_word = 16'h748f;
			12'h74a: tri_word = 16'h749f;
			12'h74b: tri_word = 16'h74af;
			12'h74c: tri_word = 16'h74bf;
			12'h74d: tri_word = 16'h74cf;
			12'h74e: tri_word = 16'h74df;
			12'h74f: tri_word = 16'h74ef;
			12'h750: tri_word = 16'h74ff;
			12'h751: tri_word = 16'h750f;
			12'h752: tri_word = 16'h751f;
			12'h753: tri_word = 16'h752f;
			12'h754: tri_word = 16'h753f;
			12'h755: tri_word = 16'h754f;
			12'h756: tri_word = 16'h755f;
			12'h757: tri_word = 16'h756f;
			12'h758: tri_word = 16'h757f;
			12'h759: tri_word = 16'h758f;
			12'h75a: tri_word = 16'h759f;
			12'h75b: tri_word = 16'h75af;
			12'h75c: tri_word = 16'h75bf;
			12'h75d: tri_word = 16'h75cf;
			12'h75e: tri_word = 16'h75df;
			12'h75f: tri_word = 16'h75ef;
			12'h760: tri_word = 16'h75ff;
			12'h761: tri_word = 16'h760f;
			12'h762: tri_word = 16'h761f;
			12'h763: tri_word = 16'h762f;
			12'h764: tri_word = 16'h763f;
			12'h765: tri_word = 16'h764f;
			12'h766: tri_word = 16'h765f;
			12'h767: tri_word = 16'h766f;
			12'h768: tri_word = 16'h767f;
			12'h769: tri_word = 16'h768f;
			12'h76a: tri_word = 16'h769f;
			12'h76b: tri_word = 16'h76af;
			12'h76c: tri_word = 16'h76bf;
			12'h76d: tri_word = 16'h76cf;
			12'h76e: tri_word = 16'h76df;
			12'h76f: tri_word = 16'h76ef;
			12'h770: tri_word = 16'h76ff;
			12'h771: tri_word = 16'h770f;
			12'h772: tri_word = 16'h771f;
			12'h773: tri_word = 16'h772f;
			12'h774: tri_word = 16'h773f;
			12'h775: tri_word = 16'h774f;
			12'h776: tri_word = 16'h775f;
			12'h777: tri_word = 16'h776f;
			12'h778: tri_word = 16'h777f;
			12'h779: tri_word = 16'h778f;
			12'h77a: tri_word = 16'h779f;
			12'h77b: tri_word = 16'h77af;
			12'h77c: tri_word = 16'h77bf;
			12'h77d: tri_word = 16'h77cf;
			12'h77e: tri_word = 16'h77df;
			12'h77f: tri_word = 16'h77ef;
			12'h780: tri_word = 16'h77ff;
			12'h781: tri_word = 16'h780f;
			12'h782: tri_word = 16'h781f;
			12'h783: tri_word = 16'h782f;
			12'h784: tri_word = 16'h783f;
			12'h785: tri_word = 16'h784f;
			12'h786: tri_word = 16'h785f;
			12'h787: tri_word = 16'h786f;
			12'h788: tri_word = 16'h787f;
			12'h789: tri_word = 16'h788f;
			12'h78a: tri_word = 16'h789f;
			12'h78b: tri_word = 16'h78af;
			12'h78c: tri_word = 16'h78bf;
			12'h78d: tri_word = 16'h78cf;
			12'h78e: tri_word = 16'h78df;
			12'h78f: tri_word = 16'h78ef;
			12'h790: tri_word = 16'h78ff;
			12'h791: tri_word = 16'h790f;
			12'h792: tri_word = 16'h791f;
			12'h793: tri_word = 16'h792f;
			12'h794: tri_word = 16'h793f;
			12'h795: tri_word = 16'h794f;
			12'h796: tri_word = 16'h795f;
			12'h797: tri_word = 16'h796f;
			12'h798: tri_word = 16'h797f;
			12'h799: tri_word = 16'h798f;
			12'h79a: tri_word = 16'h799f;
			12'h79b: tri_word = 16'h79af;
			12'h79c: tri_word = 16'h79bf;
			12'h79d: tri_word = 16'h79cf;
			12'h79e: tri_word = 16'h79df;
			12'h79f: tri_word = 16'h79ef;
			12'h7a0: tri_word = 16'h79ff;
			12'h7a1: tri_word = 16'h7a0f;
			12'h7a2: tri_word = 16'h7a1f;
			12'h7a3: tri_word = 16'h7a2f;
			12'h7a4: tri_word = 16'h7a3f;
			12'h7a5: tri_word = 16'h7a4f;
			12'h7a6: tri_word = 16'h7a5f;
			12'h7a7: tri_word = 16'h7a6f;
			12'h7a8: tri_word = 16'h7a7f;
			12'h7a9: tri_word = 16'h7a8f;
			12'h7aa: tri_word = 16'h7a9f;
			12'h7ab: tri_word = 16'h7aaf;
			12'h7ac: tri_word = 16'h7abf;
			12'h7ad: tri_word = 16'h7acf;
			12'h7ae: tri_word = 16'h7adf;
			12'h7af: tri_word = 16'h7aef;
			12'h7b0: tri_word = 16'h7aff;
			12'h7b1: tri_word = 16'h7b0f;
			12'h7b2: tri_word = 16'h7b1f;
			12'h7b3: tri_word = 16'h7b2f;
			12'h7b4: tri_word = 16'h7b3f;
			12'h7b5: tri_word = 16'h7b4f;
			12'h7b6: tri_word = 16'h7b5f;
			12'h7b7: tri_word = 16'h7b6f;
			12'h7b8: tri_word = 16'h7b7f;
			12'h7b9: tri_word = 16'h7b8f;
			12'h7ba: tri_word = 16'h7b9f;
			12'h7bb: tri_word = 16'h7baf;
			12'h7bc: tri_word = 16'h7bbf;
			12'h7bd: tri_word = 16'h7bcf;
			12'h7be: tri_word = 16'h7bdf;
			12'h7bf: tri_word = 16'h7bef;
			12'h7c0: tri_word = 16'h7bff;
			12'h7c1: tri_word = 16'h7c0f;
			12'h7c2: tri_word = 16'h7c1f;
			12'h7c3: tri_word = 16'h7c2f;
			12'h7c4: tri_word = 16'h7c3f;
			12'h7c5: tri_word = 16'h7c4f;
			12'h7c6: tri_word = 16'h7c5f;
			12'h7c7: tri_word = 16'h7c6f;
			12'h7c8: tri_word = 16'h7c7f;
			12'h7c9: tri_word = 16'h7c8f;
			12'h7ca: tri_word = 16'h7c9f;
			12'h7cb: tri_word = 16'h7caf;
			12'h7cc: tri_word = 16'h7cbf;
			12'h7cd: tri_word = 16'h7ccf;
			12'h7ce: tri_word = 16'h7cdf;
			12'h7cf: tri_word = 16'h7cef;
			12'h7d0: tri_word = 16'h7cff;
			12'h7d1: tri_word = 16'h7d0f;
			12'h7d2: tri_word = 16'h7d1f;
			12'h7d3: tri_word = 16'h7d2f;
			12'h7d4: tri_word = 16'h7d3f;
			12'h7d5: tri_word = 16'h7d4f;
			12'h7d6: tri_word = 16'h7d5f;
			12'h7d7: tri_word = 16'h7d6f;
			12'h7d8: tri_word = 16'h7d7f;
			12'h7d9: tri_word = 16'h7d8f;
			12'h7da: tri_word = 16'h7d9f;
			12'h7db: tri_word = 16'h7daf;
			12'h7dc: tri_word = 16'h7dbf;
			12'h7dd: tri_word = 16'h7dcf;
			12'h7de: tri_word = 16'h7ddf;
			12'h7df: tri_word = 16'h7def;
			12'h7e0: tri_word = 16'h7dff;
			12'h7e1: tri_word = 16'h7e0f;
			12'h7e2: tri_word = 16'h7e1f;
			12'h7e3: tri_word = 16'h7e2f;
			12'h7e4: tri_word = 16'h7e3f;
			12'h7e5: tri_word = 16'h7e4f;
			12'h7e6: tri_word = 16'h7e5f;
			12'h7e7: tri_word = 16'h7e6f;
			12'h7e8: tri_word = 16'h7e7f;
			12'h7e9: tri_word = 16'h7e8f;
			12'h7ea: tri_word = 16'h7e9f;
			12'h7eb: tri_word = 16'h7eaf;
			12'h7ec: tri_word = 16'h7ebf;
			12'h7ed: tri_word = 16'h7ecf;
			12'h7ee: tri_word = 16'h7edf;
			12'h7ef: tri_word = 16'h7eef;
			12'h7f0: tri_word = 16'h7eff;
			12'h7f1: tri_word = 16'h7f0e;
			12'h7f2: tri_word = 16'h7f1e;
			12'h7f3: tri_word = 16'h7f2e;
			12'h7f4: tri_word = 16'h7f3e;
			12'h7f5: tri_word = 16'h7f4e;
			12'h7f6: tri_word = 16'h7f5e;
			12'h7f7: tri_word = 16'h7f6e;
			12'h7f8: tri_word = 16'h7f7e;
			12'h7f9: tri_word = 16'h7f8e;
			12'h7fa: tri_word = 16'h7f9e;
			12'h7fb: tri_word = 16'h7fae;
			12'h7fc: tri_word = 16'h7fbe;
			12'h7fd: tri_word = 16'h7fce;
			12'h7fe: tri_word = 16'h7fde;
			12'h7ff: tri_word = 16'h7fee;
			12'h800: tri_word = 16'h7fff;
			12'h801: tri_word = 16'h7fef;
			12'h802: tri_word = 16'h7fdf;
			12'h803: tri_word = 16'h7fcf;
			12'h804: tri_word = 16'h7fbf;
			12'h805: tri_word = 16'h7faf;
			12'h806: tri_word = 16'h7f9f;
			12'h807: tri_word = 16'h7f8f;
			12'h808: tri_word = 16'h7f7f;
			12'h809: tri_word = 16'h7f6f;
			12'h80a: tri_word = 16'h7f5f;
			12'h80b: tri_word = 16'h7f4f;
			12'h80c: tri_word = 16'h7f3f;
			12'h80d: tri_word = 16'h7f2f;
			12'h80e: tri_word = 16'h7f1f;
			12'h80f: tri_word = 16'h7f0f;
			12'h810: tri_word = 16'h7eff;
			12'h811: tri_word = 16'h7eef;
			12'h812: tri_word = 16'h7edf;
			12'h813: tri_word = 16'h7ecf;
			12'h814: tri_word = 16'h7ebf;
			12'h815: tri_word = 16'h7eaf;
			12'h816: tri_word = 16'h7e9f;
			12'h817: tri_word = 16'h7e8f;
			12'h818: tri_word = 16'h7e7f;
			12'h819: tri_word = 16'h7e6f;
			12'h81a: tri_word = 16'h7e5f;
			12'h81b: tri_word = 16'h7e4f;
			12'h81c: tri_word = 16'h7e3f;
			12'h81d: tri_word = 16'h7e2f;
			12'h81e: tri_word = 16'h7e1f;
			12'h81f: tri_word = 16'h7e0f;
			12'h820: tri_word = 16'h7dff;
			12'h821: tri_word = 16'h7def;
			12'h822: tri_word = 16'h7ddf;
			12'h823: tri_word = 16'h7dcf;
			12'h824: tri_word = 16'h7dbf;
			12'h825: tri_word = 16'h7daf;
			12'h826: tri_word = 16'h7d9f;
			12'h827: tri_word = 16'h7d8f;
			12'h828: tri_word = 16'h7d7f;
			12'h829: tri_word = 16'h7d6f;
			12'h82a: tri_word = 16'h7d5f;
			12'h82b: tri_word = 16'h7d4f;
			12'h82c: tri_word = 16'h7d3f;
			12'h82d: tri_word = 16'h7d2f;
			12'h82e: tri_word = 16'h7d1f;
			12'h82f: tri_word = 16'h7d0f;
			12'h830: tri_word = 16'h7cff;
			12'h831: tri_word = 16'h7cef;
			12'h832: tri_word = 16'h7cdf;
			12'h833: tri_word = 16'h7ccf;
			12'h834: tri_word = 16'h7cbf;
			12'h835: tri_word = 16'h7caf;
			12'h836: tri_word = 16'h7c9f;
			12'h837: tri_word = 16'h7c8f;
			12'h838: tri_word = 16'h7c7f;
			12'h839: tri_word = 16'h7c6f;
			12'h83a: tri_word = 16'h7c5f;
			12'h83b: tri_word = 16'h7c4f;
			12'h83c: tri_word = 16'h7c3f;
			12'h83d: tri_word = 16'h7c2f;
			12'h83e: tri_word = 16'h7c1f;
			12'h83f: tri_word = 16'h7c0f;
			12'h840: tri_word = 16'h7bff;
			12'h841: tri_word = 16'h7bef;
			12'h842: tri_word = 16'h7bdf;
			12'h843: tri_word = 16'h7bcf;
			12'h844: tri_word = 16'h7bbf;
			12'h845: tri_word = 16'h7baf;
			12'h846: tri_word = 16'h7b9f;
			12'h847: tri_word = 16'h7b8f;
			12'h848: tri_word = 16'h7b7f;
			12'h849: tri_word = 16'h7b6f;
			12'h84a: tri_word = 16'h7b5f;
			12'h84b: tri_word = 16'h7b4f;
			12'h84c: tri_word = 16'h7b3f;
			12'h84d: tri_word = 16'h7b2f;
			12'h84e: tri_word = 16'h7b1f;
			12'h84f: tri_word = 16'h7b0f;
			12'h850: tri_word = 16'h7aff;
			12'h851: tri_word = 16'h7aef;
			12'h852: tri_word = 16'h7adf;
			12'h853: tri_word = 16'h7acf;
			12'h854: tri_word = 16'h7abf;
			12'h855: tri_word = 16'h7aaf;
			12'h856: tri_word = 16'h7a9f;
			12'h857: tri_word = 16'h7a8f;
			12'h858: tri_word = 16'h7a7f;
			12'h859: tri_word = 16'h7a6f;
			12'h85a: tri_word = 16'h7a5f;
			12'h85b: tri_word = 16'h7a4f;
			12'h85c: tri_word = 16'h7a3f;
			12'h85d: tri_word = 16'h7a2f;
			12'h85e: tri_word = 16'h7a1f;
			12'h85f: tri_word = 16'h7a0f;
			12'h860: tri_word = 16'h79ff;
			12'h861: tri_word = 16'h79ef;
			12'h862: tri_word = 16'h79df;
			12'h863: tri_word = 16'h79cf;
			12'h864: tri_word = 16'h79bf;
			12'h865: tri_word = 16'h79af;
			12'h866: tri_word = 16'h799f;
			12'h867: tri_word = 16'h798f;
			12'h868: tri_word = 16'h797f;
			12'h869: tri_word = 16'h796f;
			12'h86a: tri_word = 16'h795f;
			12'h86b: tri_word = 16'h794f;
			12'h86c: tri_word = 16'h793f;
			12'h86d: tri_word = 16'h792f;
			12'h86e: tri_word = 16'h791f;
			12'h86f: tri_word = 16'h790f;
			12'h870: tri_word = 16'h78ff;
			12'h871: tri_word = 16'h78ef;
			12'h872: tri_word = 16'h78df;
			12'h873: tri_word = 16'h78cf;
			12'h874: tri_word = 16'h78bf;
			12'h875: tri_word = 16'h78af;
			12'h876: tri_word = 16'h789f;
			12'h877: tri_word = 16'h788f;
			12'h878: tri_word = 16'h787f;
			12'h879: tri_word = 16'h786f;
			12'h87a: tri_word = 16'h785f;
			12'h87b: tri_word = 16'h784f;
			12'h87c: tri_word = 16'h783f;
			12'h87d: tri_word = 16'h782f;
			12'h87e: tri_word = 16'h781f;
			12'h87f: tri_word = 16'h780f;
			12'h880: tri_word = 16'h77ff;
			12'h881: tri_word = 16'h77ef;
			12'h882: tri_word = 16'h77df;
			12'h883: tri_word = 16'h77cf;
			12'h884: tri_word = 16'h77bf;
			12'h885: tri_word = 16'h77af;
			12'h886: tri_word = 16'h779f;
			12'h887: tri_word = 16'h778f;
			12'h888: tri_word = 16'h777f;
			12'h889: tri_word = 16'h776f;
			12'h88a: tri_word = 16'h775f;
			12'h88b: tri_word = 16'h774f;
			12'h88c: tri_word = 16'h773f;
			12'h88d: tri_word = 16'h772f;
			12'h88e: tri_word = 16'h771f;
			12'h88f: tri_word = 16'h770f;
			12'h890: tri_word = 16'h76ff;
			12'h891: tri_word = 16'h76ef;
			12'h892: tri_word = 16'h76df;
			12'h893: tri_word = 16'h76cf;
			12'h894: tri_word = 16'h76bf;
			12'h895: tri_word = 16'h76af;
			12'h896: tri_word = 16'h769f;
			12'h897: tri_word = 16'h768f;
			12'h898: tri_word = 16'h767f;
			12'h899: tri_word = 16'h766f;
			12'h89a: tri_word = 16'h765f;
			12'h89b: tri_word = 16'h764f;
			12'h89c: tri_word = 16'h763f;
			12'h89d: tri_word = 16'h762f;
			12'h89e: tri_word = 16'h761f;
			12'h89f: tri_word = 16'h760f;
			12'h8a0: tri_word = 16'h75ff;
			12'h8a1: tri_word = 16'h75ef;
			12'h8a2: tri_word = 16'h75df;
			12'h8a3: tri_word = 16'h75cf;
			12'h8a4: tri_word = 16'h75bf;
			12'h8a5: tri_word = 16'h75af;
			12'h8a6: tri_word = 16'h759f;
			12'h8a7: tri_word = 16'h758f;
			12'h8a8: tri_word = 16'h757f;
			12'h8a9: tri_word = 16'h756f;
			12'h8aa: tri_word = 16'h755f;
			12'h8ab: tri_word = 16'h754f;
			12'h8ac: tri_word = 16'h753f;
			12'h8ad: tri_word = 16'h752f;
			12'h8ae: tri_word = 16'h751f;
			12'h8af: tri_word = 16'h750f;
			12'h8b0: tri_word = 16'h74ff;
			12'h8b1: tri_word = 16'h74ef;
			12'h8b2: tri_word = 16'h74df;
			12'h8b3: tri_word = 16'h74cf;
			12'h8b4: tri_word = 16'h74bf;
			12'h8b5: tri_word = 16'h74af;
			12'h8b6: tri_word = 16'h749f;
			12'h8b7: tri_word = 16'h748f;
			12'h8b8: tri_word = 16'h747f;
			12'h8b9: tri_word = 16'h746f;
			12'h8ba: tri_word = 16'h745f;
			12'h8bb: tri_word = 16'h744f;
			12'h8bc: tri_word = 16'h743f;
			12'h8bd: tri_word = 16'h742f;
			12'h8be: tri_word = 16'h741f;
			12'h8bf: tri_word = 16'h740f;
			12'h8c0: tri_word = 16'h73ff;
			12'h8c1: tri_word = 16'h73ef;
			12'h8c2: tri_word = 16'h73df;
			12'h8c3: tri_word = 16'h73cf;
			12'h8c4: tri_word = 16'h73bf;
			12'h8c5: tri_word = 16'h73af;
			12'h8c6: tri_word = 16'h739f;
			12'h8c7: tri_word = 16'h738f;
			12'h8c8: tri_word = 16'h737f;
			12'h8c9: tri_word = 16'h736f;
			12'h8ca: tri_word = 16'h735f;
			12'h8cb: tri_word = 16'h734f;
			12'h8cc: tri_word = 16'h733f;
			12'h8cd: tri_word = 16'h732f;
			12'h8ce: tri_word = 16'h731f;
			12'h8cf: tri_word = 16'h730f;
			12'h8d0: tri_word = 16'h72ff;
			12'h8d1: tri_word = 16'h72ef;
			12'h8d2: tri_word = 16'h72df;
			12'h8d3: tri_word = 16'h72cf;
			12'h8d4: tri_word = 16'h72bf;
			12'h8d5: tri_word = 16'h72af;
			12'h8d6: tri_word = 16'h729f;
			12'h8d7: tri_word = 16'h728f;
			12'h8d8: tri_word = 16'h727f;
			12'h8d9: tri_word = 16'h726f;
			12'h8da: tri_word = 16'h725f;
			12'h8db: tri_word = 16'h724f;
			12'h8dc: tri_word = 16'h723f;
			12'h8dd: tri_word = 16'h722f;
			12'h8de: tri_word = 16'h721f;
			12'h8df: tri_word = 16'h720f;
			12'h8e0: tri_word = 16'h71ff;
			12'h8e1: tri_word = 16'h71ef;
			12'h8e2: tri_word = 16'h71df;
			12'h8e3: tri_word = 16'h71cf;
			12'h8e4: tri_word = 16'h71bf;
			12'h8e5: tri_word = 16'h71af;
			12'h8e6: tri_word = 16'h719f;
			12'h8e7: tri_word = 16'h718f;
			12'h8e8: tri_word = 16'h717f;
			12'h8e9: tri_word = 16'h716f;
			12'h8ea: tri_word = 16'h715f;
			12'h8eb: tri_word = 16'h714f;
			12'h8ec: tri_word = 16'h713f;
			12'h8ed: tri_word = 16'h712f;
			12'h8ee: tri_word = 16'h711f;
			12'h8ef: tri_word = 16'h710f;
			12'h8f0: tri_word = 16'h70ff;
			12'h8f1: tri_word = 16'h70ef;
			12'h8f2: tri_word = 16'h70df;
			12'h8f3: tri_word = 16'h70cf;
			12'h8f4: tri_word = 16'h70bf;
			12'h8f5: tri_word = 16'h70af;
			12'h8f6: tri_word = 16'h709f;
			12'h8f7: tri_word = 16'h708f;
			12'h8f8: tri_word = 16'h707f;
			12'h8f9: tri_word = 16'h706f;
			12'h8fa: tri_word = 16'h705f;
			12'h8fb: tri_word = 16'h704f;
			12'h8fc: tri_word = 16'h703f;
			12'h8fd: tri_word = 16'h702f;
			12'h8fe: tri_word = 16'h701f;
			12'h8ff: tri_word = 16'h700f;
			12'h900: tri_word = 16'h6fff;
			12'h901: tri_word = 16'h6fef;
			12'h902: tri_word = 16'h6fdf;
			12'h903: tri_word = 16'h6fcf;
			12'h904: tri_word = 16'h6fbf;
			12'h905: tri_word = 16'h6faf;
			12'h906: tri_word = 16'h6f9f;
			12'h907: tri_word = 16'h6f8f;
			12'h908: tri_word = 16'h6f7f;
			12'h909: tri_word = 16'h6f6f;
			12'h90a: tri_word = 16'h6f5f;
			12'h90b: tri_word = 16'h6f4f;
			12'h90c: tri_word = 16'h6f3f;
			12'h90d: tri_word = 16'h6f2f;
			12'h90e: tri_word = 16'h6f1f;
			12'h90f: tri_word = 16'h6f0f;
			12'h910: tri_word = 16'h6eff;
			12'h911: tri_word = 16'h6eef;
			12'h912: tri_word = 16'h6edf;
			12'h913: tri_word = 16'h6ecf;
			12'h914: tri_word = 16'h6ebf;
			12'h915: tri_word = 16'h6eaf;
			12'h916: tri_word = 16'h6e9f;
			12'h917: tri_word = 16'h6e8f;
			12'h918: tri_word = 16'h6e7f;
			12'h919: tri_word = 16'h6e6f;
			12'h91a: tri_word = 16'h6e5f;
			12'h91b: tri_word = 16'h6e4f;
			12'h91c: tri_word = 16'h6e3f;
			12'h91d: tri_word = 16'h6e2f;
			12'h91e: tri_word = 16'h6e1f;
			12'h91f: tri_word = 16'h6e0f;
			12'h920: tri_word = 16'h6dff;
			12'h921: tri_word = 16'h6def;
			12'h922: tri_word = 16'h6ddf;
			12'h923: tri_word = 16'h6dcf;
			12'h924: tri_word = 16'h6dbf;
			12'h925: tri_word = 16'h6daf;
			12'h926: tri_word = 16'h6d9f;
			12'h927: tri_word = 16'h6d8f;
			12'h928: tri_word = 16'h6d7f;
			12'h929: tri_word = 16'h6d6f;
			12'h92a: tri_word = 16'h6d5f;
			12'h92b: tri_word = 16'h6d4f;
			12'h92c: tri_word = 16'h6d3f;
			12'h92d: tri_word = 16'h6d2f;
			12'h92e: tri_word = 16'h6d1f;
			12'h92f: tri_word = 16'h6d0f;
			12'h930: tri_word = 16'h6cff;
			12'h931: tri_word = 16'h6cef;
			12'h932: tri_word = 16'h6cdf;
			12'h933: tri_word = 16'h6ccf;
			12'h934: tri_word = 16'h6cbf;
			12'h935: tri_word = 16'h6caf;
			12'h936: tri_word = 16'h6c9f;
			12'h937: tri_word = 16'h6c8f;
			12'h938: tri_word = 16'h6c7f;
			12'h939: tri_word = 16'h6c6f;
			12'h93a: tri_word = 16'h6c5f;
			12'h93b: tri_word = 16'h6c4f;
			12'h93c: tri_word = 16'h6c3f;
			12'h93d: tri_word = 16'h6c2f;
			12'h93e: tri_word = 16'h6c1f;
			12'h93f: tri_word = 16'h6c0f;
			12'h940: tri_word = 16'h6bff;
			12'h941: tri_word = 16'h6bef;
			12'h942: tri_word = 16'h6bdf;
			12'h943: tri_word = 16'h6bcf;
			12'h944: tri_word = 16'h6bbf;
			12'h945: tri_word = 16'h6baf;
			12'h946: tri_word = 16'h6b9f;
			12'h947: tri_word = 16'h6b8f;
			12'h948: tri_word = 16'h6b7f;
			12'h949: tri_word = 16'h6b6f;
			12'h94a: tri_word = 16'h6b5f;
			12'h94b: tri_word = 16'h6b4f;
			12'h94c: tri_word = 16'h6b3f;
			12'h94d: tri_word = 16'h6b2f;
			12'h94e: tri_word = 16'h6b1f;
			12'h94f: tri_word = 16'h6b0f;
			12'h950: tri_word = 16'h6aff;
			12'h951: tri_word = 16'h6aef;
			12'h952: tri_word = 16'h6adf;
			12'h953: tri_word = 16'h6acf;
			12'h954: tri_word = 16'h6abf;
			12'h955: tri_word = 16'h6aaf;
			12'h956: tri_word = 16'h6a9f;
			12'h957: tri_word = 16'h6a8f;
			12'h958: tri_word = 16'h6a7f;
			12'h959: tri_word = 16'h6a6f;
			12'h95a: tri_word = 16'h6a5f;
			12'h95b: tri_word = 16'h6a4f;
			12'h95c: tri_word = 16'h6a3f;
			12'h95d: tri_word = 16'h6a2f;
			12'h95e: tri_word = 16'h6a1f;
			12'h95f: tri_word = 16'h6a0f;
			12'h960: tri_word = 16'h69ff;
			12'h961: tri_word = 16'h69ef;
			12'h962: tri_word = 16'h69df;
			12'h963: tri_word = 16'h69cf;
			12'h964: tri_word = 16'h69bf;
			12'h965: tri_word = 16'h69af;
			12'h966: tri_word = 16'h699f;
			12'h967: tri_word = 16'h698f;
			12'h968: tri_word = 16'h697f;
			12'h969: tri_word = 16'h696f;
			12'h96a: tri_word = 16'h695f;
			12'h96b: tri_word = 16'h694f;
			12'h96c: tri_word = 16'h693f;
			12'h96d: tri_word = 16'h692f;
			12'h96e: tri_word = 16'h691f;
			12'h96f: tri_word = 16'h690f;
			12'h970: tri_word = 16'h68ff;
			12'h971: tri_word = 16'h68ef;
			12'h972: tri_word = 16'h68df;
			12'h973: tri_word = 16'h68cf;
			12'h974: tri_word = 16'h68bf;
			12'h975: tri_word = 16'h68af;
			12'h976: tri_word = 16'h689f;
			12'h977: tri_word = 16'h688f;
			12'h978: tri_word = 16'h687f;
			12'h979: tri_word = 16'h686f;
			12'h97a: tri_word = 16'h685f;
			12'h97b: tri_word = 16'h684f;
			12'h97c: tri_word = 16'h683f;
			12'h97d: tri_word = 16'h682f;
			12'h97e: tri_word = 16'h681f;
			12'h97f: tri_word = 16'h680f;
			12'h980: tri_word = 16'h67ff;
			12'h981: tri_word = 16'h67ef;
			12'h982: tri_word = 16'h67df;
			12'h983: tri_word = 16'h67cf;
			12'h984: tri_word = 16'h67bf;
			12'h985: tri_word = 16'h67af;
			12'h986: tri_word = 16'h679f;
			12'h987: tri_word = 16'h678f;
			12'h988: tri_word = 16'h677f;
			12'h989: tri_word = 16'h676f;
			12'h98a: tri_word = 16'h675f;
			12'h98b: tri_word = 16'h674f;
			12'h98c: tri_word = 16'h673f;
			12'h98d: tri_word = 16'h672f;
			12'h98e: tri_word = 16'h671f;
			12'h98f: tri_word = 16'h670f;
			12'h990: tri_word = 16'h66ff;
			12'h991: tri_word = 16'h66ef;
			12'h992: tri_word = 16'h66df;
			12'h993: tri_word = 16'h66cf;
			12'h994: tri_word = 16'h66bf;
			12'h995: tri_word = 16'h66af;
			12'h996: tri_word = 16'h669f;
			12'h997: tri_word = 16'h668f;
			12'h998: tri_word = 16'h667f;
			12'h999: tri_word = 16'h666f;
			12'h99a: tri_word = 16'h665f;
			12'h99b: tri_word = 16'h664f;
			12'h99c: tri_word = 16'h663f;
			12'h99d: tri_word = 16'h662f;
			12'h99e: tri_word = 16'h661f;
			12'h99f: tri_word = 16'h660f;
			12'h9a0: tri_word = 16'h65ff;
			12'h9a1: tri_word = 16'h65ef;
			12'h9a2: tri_word = 16'h65df;
			12'h9a3: tri_word = 16'h65cf;
			12'h9a4: tri_word = 16'h65bf;
			12'h9a5: tri_word = 16'h65af;
			12'h9a6: tri_word = 16'h659f;
			12'h9a7: tri_word = 16'h658f;
			12'h9a8: tri_word = 16'h657f;
			12'h9a9: tri_word = 16'h656f;
			12'h9aa: tri_word = 16'h655f;
			12'h9ab: tri_word = 16'h654f;
			12'h9ac: tri_word = 16'h653f;
			12'h9ad: tri_word = 16'h652f;
			12'h9ae: tri_word = 16'h651f;
			12'h9af: tri_word = 16'h650f;
			12'h9b0: tri_word = 16'h64ff;
			12'h9b1: tri_word = 16'h64ef;
			12'h9b2: tri_word = 16'h64df;
			12'h9b3: tri_word = 16'h64cf;
			12'h9b4: tri_word = 16'h64bf;
			12'h9b5: tri_word = 16'h64af;
			12'h9b6: tri_word = 16'h649f;
			12'h9b7: tri_word = 16'h648f;
			12'h9b8: tri_word = 16'h647f;
			12'h9b9: tri_word = 16'h646f;
			12'h9ba: tri_word = 16'h645f;
			12'h9bb: tri_word = 16'h644f;
			12'h9bc: tri_word = 16'h643f;
			12'h9bd: tri_word = 16'h642f;
			12'h9be: tri_word = 16'h641f;
			12'h9bf: tri_word = 16'h640f;
			12'h9c0: tri_word = 16'h63ff;
			12'h9c1: tri_word = 16'h63ef;
			12'h9c2: tri_word = 16'h63df;
			12'h9c3: tri_word = 16'h63cf;
			12'h9c4: tri_word = 16'h63bf;
			12'h9c5: tri_word = 16'h63af;
			12'h9c6: tri_word = 16'h639f;
			12'h9c7: tri_word = 16'h638f;
			12'h9c8: tri_word = 16'h637f;
			12'h9c9: tri_word = 16'h636f;
			12'h9ca: tri_word = 16'h635f;
			12'h9cb: tri_word = 16'h634f;
			12'h9cc: tri_word = 16'h633f;
			12'h9cd: tri_word = 16'h632f;
			12'h9ce: tri_word = 16'h631f;
			12'h9cf: tri_word = 16'h630f;
			12'h9d0: tri_word = 16'h62ff;
			12'h9d1: tri_word = 16'h62ef;
			12'h9d2: tri_word = 16'h62df;
			12'h9d3: tri_word = 16'h62cf;
			12'h9d4: tri_word = 16'h62bf;
			12'h9d5: tri_word = 16'h62af;
			12'h9d6: tri_word = 16'h629f;
			12'h9d7: tri_word = 16'h628f;
			12'h9d8: tri_word = 16'h627f;
			12'h9d9: tri_word = 16'h626f;
			12'h9da: tri_word = 16'h625f;
			12'h9db: tri_word = 16'h624f;
			12'h9dc: tri_word = 16'h623f;
			12'h9dd: tri_word = 16'h622f;
			12'h9de: tri_word = 16'h621f;
			12'h9df: tri_word = 16'h620f;
			12'h9e0: tri_word = 16'h61ff;
			12'h9e1: tri_word = 16'h61ef;
			12'h9e2: tri_word = 16'h61df;
			12'h9e3: tri_word = 16'h61cf;
			12'h9e4: tri_word = 16'h61bf;
			12'h9e5: tri_word = 16'h61af;
			12'h9e6: tri_word = 16'h619f;
			12'h9e7: tri_word = 16'h618f;
			12'h9e8: tri_word = 16'h617f;
			12'h9e9: tri_word = 16'h616f;
			12'h9ea: tri_word = 16'h615f;
			12'h9eb: tri_word = 16'h614f;
			12'h9ec: tri_word = 16'h613f;
			12'h9ed: tri_word = 16'h612f;
			12'h9ee: tri_word = 16'h611f;
			12'h9ef: tri_word = 16'h610f;
			12'h9f0: tri_word = 16'h60ff;
			12'h9f1: tri_word = 16'h60ef;
			12'h9f2: tri_word = 16'h60df;
			12'h9f3: tri_word = 16'h60cf;
			12'h9f4: tri_word = 16'h60bf;
			12'h9f5: tri_word = 16'h60af;
			12'h9f6: tri_word = 16'h609f;
			12'h9f7: tri_word = 16'h608f;
			12'h9f8: tri_word = 16'h607f;
			12'h9f9: tri_word = 16'h606f;
			12'h9fa: tri_word = 16'h605f;
			12'h9fb: tri_word = 16'h604f;
			12'h9fc: tri_word = 16'h603f;
			12'h9fd: tri_word = 16'h602f;
			12'h9fe: tri_word = 16'h601f;
			12'h9ff: tri_word = 16'h600f;
			12'ha00: tri_word = 16'h5fff;
			12'ha01: tri_word = 16'h5fef;
			12'ha02: tri_word = 16'h5fdf;
			12'ha03: tri_word = 16'h5fcf;
			12'ha04: tri_word = 16'h5fbf;
			12'ha05: tri_word = 16'h5faf;
			12'ha06: tri_word = 16'h5f9f;
			12'ha07: tri_word = 16'h5f8f;
			12'ha08: tri_word = 16'h5f7f;
			12'ha09: tri_word = 16'h5f6f;
			12'ha0a: tri_word = 16'h5f5f;
			12'ha0b: tri_word = 16'h5f4f;
			12'ha0c: tri_word = 16'h5f3f;
			12'ha0d: tri_word = 16'h5f2f;
			12'ha0e: tri_word = 16'h5f1f;
			12'ha0f: tri_word = 16'h5f0f;
			12'ha10: tri_word = 16'h5eff;
			12'ha11: tri_word = 16'h5eef;
			12'ha12: tri_word = 16'h5edf;
			12'ha13: tri_word = 16'h5ecf;
			12'ha14: tri_word = 16'h5ebf;
			12'ha15: tri_word = 16'h5eaf;
			12'ha16: tri_word = 16'h5e9f;
			12'ha17: tri_word = 16'h5e8f;
			12'ha18: tri_word = 16'h5e7f;
			12'ha19: tri_word = 16'h5e6f;
			12'ha1a: tri_word = 16'h5e5f;
			12'ha1b: tri_word = 16'h5e4f;
			12'ha1c: tri_word = 16'h5e3f;
			12'ha1d: tri_word = 16'h5e2f;
			12'ha1e: tri_word = 16'h5e1f;
			12'ha1f: tri_word = 16'h5e0f;
			12'ha20: tri_word = 16'h5dff;
			12'ha21: tri_word = 16'h5def;
			12'ha22: tri_word = 16'h5ddf;
			12'ha23: tri_word = 16'h5dcf;
			12'ha24: tri_word = 16'h5dbf;
			12'ha25: tri_word = 16'h5daf;
			12'ha26: tri_word = 16'h5d9f;
			12'ha27: tri_word = 16'h5d8f;
			12'ha28: tri_word = 16'h5d7f;
			12'ha29: tri_word = 16'h5d6f;
			12'ha2a: tri_word = 16'h5d5f;
			12'ha2b: tri_word = 16'h5d4f;
			12'ha2c: tri_word = 16'h5d3f;
			12'ha2d: tri_word = 16'h5d2f;
			12'ha2e: tri_word = 16'h5d1f;
			12'ha2f: tri_word = 16'h5d0f;
			12'ha30: tri_word = 16'h5cff;
			12'ha31: tri_word = 16'h5cef;
			12'ha32: tri_word = 16'h5cdf;
			12'ha33: tri_word = 16'h5ccf;
			12'ha34: tri_word = 16'h5cbf;
			12'ha35: tri_word = 16'h5caf;
			12'ha36: tri_word = 16'h5c9f;
			12'ha37: tri_word = 16'h5c8f;
			12'ha38: tri_word = 16'h5c7f;
			12'ha39: tri_word = 16'h5c6f;
			12'ha3a: tri_word = 16'h5c5f;
			12'ha3b: tri_word = 16'h5c4f;
			12'ha3c: tri_word = 16'h5c3f;
			12'ha3d: tri_word = 16'h5c2f;
			12'ha3e: tri_word = 16'h5c1f;
			12'ha3f: tri_word = 16'h5c0f;
			12'ha40: tri_word = 16'h5bff;
			12'ha41: tri_word = 16'h5bef;
			12'ha42: tri_word = 16'h5bdf;
			12'ha43: tri_word = 16'h5bcf;
			12'ha44: tri_word = 16'h5bbf;
			12'ha45: tri_word = 16'h5baf;
			12'ha46: tri_word = 16'h5b9f;
			12'ha47: tri_word = 16'h5b8f;
			12'ha48: tri_word = 16'h5b7f;
			12'ha49: tri_word = 16'h5b6f;
			12'ha4a: tri_word = 16'h5b5f;
			12'ha4b: tri_word = 16'h5b4f;
			12'ha4c: tri_word = 16'h5b3f;
			12'ha4d: tri_word = 16'h5b2f;
			12'ha4e: tri_word = 16'h5b1f;
			12'ha4f: tri_word = 16'h5b0f;
			12'ha50: tri_word = 16'h5aff;
			12'ha51: tri_word = 16'h5aef;
			12'ha52: tri_word = 16'h5adf;
			12'ha53: tri_word = 16'h5acf;
			12'ha54: tri_word = 16'h5abf;
			12'ha55: tri_word = 16'h5aaf;
			12'ha56: tri_word = 16'h5a9f;
			12'ha57: tri_word = 16'h5a8f;
			12'ha58: tri_word = 16'h5a7f;
			12'ha59: tri_word = 16'h5a6f;
			12'ha5a: tri_word = 16'h5a5f;
			12'ha5b: tri_word = 16'h5a4f;
			12'ha5c: tri_word = 16'h5a3f;
			12'ha5d: tri_word = 16'h5a2f;
			12'ha5e: tri_word = 16'h5a1f;
			12'ha5f: tri_word = 16'h5a0f;
			12'ha60: tri_word = 16'h59ff;
			12'ha61: tri_word = 16'h59ef;
			12'ha62: tri_word = 16'h59df;
			12'ha63: tri_word = 16'h59cf;
			12'ha64: tri_word = 16'h59bf;
			12'ha65: tri_word = 16'h59af;
			12'ha66: tri_word = 16'h599f;
			12'ha67: tri_word = 16'h598f;
			12'ha68: tri_word = 16'h597f;
			12'ha69: tri_word = 16'h596f;
			12'ha6a: tri_word = 16'h595f;
			12'ha6b: tri_word = 16'h594f;
			12'ha6c: tri_word = 16'h593f;
			12'ha6d: tri_word = 16'h592f;
			12'ha6e: tri_word = 16'h591f;
			12'ha6f: tri_word = 16'h590f;
			12'ha70: tri_word = 16'h58ff;
			12'ha71: tri_word = 16'h58ef;
			12'ha72: tri_word = 16'h58df;
			12'ha73: tri_word = 16'h58cf;
			12'ha74: tri_word = 16'h58bf;
			12'ha75: tri_word = 16'h58af;
			12'ha76: tri_word = 16'h589f;
			12'ha77: tri_word = 16'h588f;
			12'ha78: tri_word = 16'h587f;
			12'ha79: tri_word = 16'h586f;
			12'ha7a: tri_word = 16'h585f;
			12'ha7b: tri_word = 16'h584f;
			12'ha7c: tri_word = 16'h583f;
			12'ha7d: tri_word = 16'h582f;
			12'ha7e: tri_word = 16'h581f;
			12'ha7f: tri_word = 16'h580f;
			12'ha80: tri_word = 16'h57ff;
			12'ha81: tri_word = 16'h57ef;
			12'ha82: tri_word = 16'h57df;
			12'ha83: tri_word = 16'h57cf;
			12'ha84: tri_word = 16'h57bf;
			12'ha85: tri_word = 16'h57af;
			12'ha86: tri_word = 16'h579f;
			12'ha87: tri_word = 16'h578f;
			12'ha88: tri_word = 16'h577f;
			12'ha89: tri_word = 16'h576f;
			12'ha8a: tri_word = 16'h575f;
			12'ha8b: tri_word = 16'h574f;
			12'ha8c: tri_word = 16'h573f;
			12'ha8d: tri_word = 16'h572f;
			12'ha8e: tri_word = 16'h571f;
			12'ha8f: tri_word = 16'h570f;
			12'ha90: tri_word = 16'h56ff;
			12'ha91: tri_word = 16'h56ef;
			12'ha92: tri_word = 16'h56df;
			12'ha93: tri_word = 16'h56cf;
			12'ha94: tri_word = 16'h56bf;
			12'ha95: tri_word = 16'h56af;
			12'ha96: tri_word = 16'h569f;
			12'ha97: tri_word = 16'h568f;
			12'ha98: tri_word = 16'h567f;
			12'ha99: tri_word = 16'h566f;
			12'ha9a: tri_word = 16'h565f;
			12'ha9b: tri_word = 16'h564f;
			12'ha9c: tri_word = 16'h563f;
			12'ha9d: tri_word = 16'h562f;
			12'ha9e: tri_word = 16'h561f;
			12'ha9f: tri_word = 16'h560f;
			12'haa0: tri_word = 16'h55ff;
			12'haa1: tri_word = 16'h55ef;
			12'haa2: tri_word = 16'h55df;
			12'haa3: tri_word = 16'h55cf;
			12'haa4: tri_word = 16'h55bf;
			12'haa5: tri_word = 16'h55af;
			12'haa6: tri_word = 16'h559f;
			12'haa7: tri_word = 16'h558f;
			12'haa8: tri_word = 16'h557f;
			12'haa9: tri_word = 16'h556f;
			12'haaa: tri_word = 16'h555f;
			12'haab: tri_word = 16'h554f;
			12'haac: tri_word = 16'h553f;
			12'haad: tri_word = 16'h552f;
			12'haae: tri_word = 16'h551f;
			12'haaf: tri_word = 16'h550f;
			12'hab0: tri_word = 16'h54ff;
			12'hab1: tri_word = 16'h54ef;
			12'hab2: tri_word = 16'h54df;
			12'hab3: tri_word = 16'h54cf;
			12'hab4: tri_word = 16'h54bf;
			12'hab5: tri_word = 16'h54af;
			12'hab6: tri_word = 16'h549f;
			12'hab7: tri_word = 16'h548f;
			12'hab8: tri_word = 16'h547f;
			12'hab9: tri_word = 16'h546f;
			12'haba: tri_word = 16'h545f;
			12'habb: tri_word = 16'h544f;
			12'habc: tri_word = 16'h543f;
			12'habd: tri_word = 16'h542f;
			12'habe: tri_word = 16'h541f;
			12'habf: tri_word = 16'h540f;
			12'hac0: tri_word = 16'h53ff;
			12'hac1: tri_word = 16'h53ef;
			12'hac2: tri_word = 16'h53df;
			12'hac3: tri_word = 16'h53cf;
			12'hac4: tri_word = 16'h53bf;
			12'hac5: tri_word = 16'h53af;
			12'hac6: tri_word = 16'h539f;
			12'hac7: tri_word = 16'h538f;
			12'hac8: tri_word = 16'h537f;
			12'hac9: tri_word = 16'h536f;
			12'haca: tri_word = 16'h535f;
			12'hacb: tri_word = 16'h534f;
			12'hacc: tri_word = 16'h533f;
			12'hacd: tri_word = 16'h532f;
			12'hace: tri_word = 16'h531f;
			12'hacf: tri_word = 16'h530f;
			12'had0: tri_word = 16'h52ff;
			12'had1: tri_word = 16'h52ef;
			12'had2: tri_word = 16'h52df;
			12'had3: tri_word = 16'h52cf;
			12'had4: tri_word = 16'h52bf;
			12'had5: tri_word = 16'h52af;
			12'had6: tri_word = 16'h529f;
			12'had7: tri_word = 16'h528f;
			12'had8: tri_word = 16'h527f;
			12'had9: tri_word = 16'h526f;
			12'hada: tri_word = 16'h525f;
			12'hadb: tri_word = 16'h524f;
			12'hadc: tri_word = 16'h523f;
			12'hadd: tri_word = 16'h522f;
			12'hade: tri_word = 16'h521f;
			12'hadf: tri_word = 16'h520f;
			12'hae0: tri_word = 16'h51ff;
			12'hae1: tri_word = 16'h51ef;
			12'hae2: tri_word = 16'h51df;
			12'hae3: tri_word = 16'h51cf;
			12'hae4: tri_word = 16'h51bf;
			12'hae5: tri_word = 16'h51af;
			12'hae6: tri_word = 16'h519f;
			12'hae7: tri_word = 16'h518f;
			12'hae8: tri_word = 16'h517f;
			12'hae9: tri_word = 16'h516f;
			12'haea: tri_word = 16'h515f;
			12'haeb: tri_word = 16'h514f;
			12'haec: tri_word = 16'h513f;
			12'haed: tri_word = 16'h512f;
			12'haee: tri_word = 16'h511f;
			12'haef: tri_word = 16'h510f;
			12'haf0: tri_word = 16'h50ff;
			12'haf1: tri_word = 16'h50ef;
			12'haf2: tri_word = 16'h50df;
			12'haf3: tri_word = 16'h50cf;
			12'haf4: tri_word = 16'h50bf;
			12'haf5: tri_word = 16'h50af;
			12'haf6: tri_word = 16'h509f;
			12'haf7: tri_word = 16'h508f;
			12'haf8: tri_word = 16'h507f;
			12'haf9: tri_word = 16'h506f;
			12'hafa: tri_word = 16'h505f;
			12'hafb: tri_word = 16'h504f;
			12'hafc: tri_word = 16'h503f;
			12'hafd: tri_word = 16'h502f;
			12'hafe: tri_word = 16'h501f;
			12'haff: tri_word = 16'h500f;
			12'hb00: tri_word = 16'h4fff;
			12'hb01: tri_word = 16'h4fef;
			12'hb02: tri_word = 16'h4fdf;
			12'hb03: tri_word = 16'h4fcf;
			12'hb04: tri_word = 16'h4fbf;
			12'hb05: tri_word = 16'h4faf;
			12'hb06: tri_word = 16'h4f9f;
			12'hb07: tri_word = 16'h4f8f;
			12'hb08: tri_word = 16'h4f7f;
			12'hb09: tri_word = 16'h4f6f;
			12'hb0a: tri_word = 16'h4f5f;
			12'hb0b: tri_word = 16'h4f4f;
			12'hb0c: tri_word = 16'h4f3f;
			12'hb0d: tri_word = 16'h4f2f;
			12'hb0e: tri_word = 16'h4f1f;
			12'hb0f: tri_word = 16'h4f0f;
			12'hb10: tri_word = 16'h4eff;
			12'hb11: tri_word = 16'h4eef;
			12'hb12: tri_word = 16'h4edf;
			12'hb13: tri_word = 16'h4ecf;
			12'hb14: tri_word = 16'h4ebf;
			12'hb15: tri_word = 16'h4eaf;
			12'hb16: tri_word = 16'h4e9f;
			12'hb17: tri_word = 16'h4e8f;
			12'hb18: tri_word = 16'h4e7f;
			12'hb19: tri_word = 16'h4e6f;
			12'hb1a: tri_word = 16'h4e5f;
			12'hb1b: tri_word = 16'h4e4f;
			12'hb1c: tri_word = 16'h4e3f;
			12'hb1d: tri_word = 16'h4e2f;
			12'hb1e: tri_word = 16'h4e1f;
			12'hb1f: tri_word = 16'h4e0f;
			12'hb20: tri_word = 16'h4dff;
			12'hb21: tri_word = 16'h4def;
			12'hb22: tri_word = 16'h4ddf;
			12'hb23: tri_word = 16'h4dcf;
			12'hb24: tri_word = 16'h4dbf;
			12'hb25: tri_word = 16'h4daf;
			12'hb26: tri_word = 16'h4d9f;
			12'hb27: tri_word = 16'h4d8f;
			12'hb28: tri_word = 16'h4d7f;
			12'hb29: tri_word = 16'h4d6f;
			12'hb2a: tri_word = 16'h4d5f;
			12'hb2b: tri_word = 16'h4d4f;
			12'hb2c: tri_word = 16'h4d3f;
			12'hb2d: tri_word = 16'h4d2f;
			12'hb2e: tri_word = 16'h4d1f;
			12'hb2f: tri_word = 16'h4d0f;
			12'hb30: tri_word = 16'h4cff;
			12'hb31: tri_word = 16'h4cef;
			12'hb32: tri_word = 16'h4cdf;
			12'hb33: tri_word = 16'h4ccf;
			12'hb34: tri_word = 16'h4cbf;
			12'hb35: tri_word = 16'h4caf;
			12'hb36: tri_word = 16'h4c9f;
			12'hb37: tri_word = 16'h4c8f;
			12'hb38: tri_word = 16'h4c7f;
			12'hb39: tri_word = 16'h4c6f;
			12'hb3a: tri_word = 16'h4c5f;
			12'hb3b: tri_word = 16'h4c4f;
			12'hb3c: tri_word = 16'h4c3f;
			12'hb3d: tri_word = 16'h4c2f;
			12'hb3e: tri_word = 16'h4c1f;
			12'hb3f: tri_word = 16'h4c0f;
			12'hb40: tri_word = 16'h4bff;
			12'hb41: tri_word = 16'h4bef;
			12'hb42: tri_word = 16'h4bdf;
			12'hb43: tri_word = 16'h4bcf;
			12'hb44: tri_word = 16'h4bbf;
			12'hb45: tri_word = 16'h4baf;
			12'hb46: tri_word = 16'h4b9f;
			12'hb47: tri_word = 16'h4b8f;
			12'hb48: tri_word = 16'h4b7f;
			12'hb49: tri_word = 16'h4b6f;
			12'hb4a: tri_word = 16'h4b5f;
			12'hb4b: tri_word = 16'h4b4f;
			12'hb4c: tri_word = 16'h4b3f;
			12'hb4d: tri_word = 16'h4b2f;
			12'hb4e: tri_word = 16'h4b1f;
			12'hb4f: tri_word = 16'h4b0f;
			12'hb50: tri_word = 16'h4aff;
			12'hb51: tri_word = 16'h4aef;
			12'hb52: tri_word = 16'h4adf;
			12'hb53: tri_word = 16'h4acf;
			12'hb54: tri_word = 16'h4abf;
			12'hb55: tri_word = 16'h4aaf;
			12'hb56: tri_word = 16'h4a9f;
			12'hb57: tri_word = 16'h4a8f;
			12'hb58: tri_word = 16'h4a7f;
			12'hb59: tri_word = 16'h4a6f;
			12'hb5a: tri_word = 16'h4a5f;
			12'hb5b: tri_word = 16'h4a4f;
			12'hb5c: tri_word = 16'h4a3f;
			12'hb5d: tri_word = 16'h4a2f;
			12'hb5e: tri_word = 16'h4a1f;
			12'hb5f: tri_word = 16'h4a0f;
			12'hb60: tri_word = 16'h49ff;
			12'hb61: tri_word = 16'h49ef;
			12'hb62: tri_word = 16'h49df;
			12'hb63: tri_word = 16'h49cf;
			12'hb64: tri_word = 16'h49bf;
			12'hb65: tri_word = 16'h49af;
			12'hb66: tri_word = 16'h499f;
			12'hb67: tri_word = 16'h498f;
			12'hb68: tri_word = 16'h497f;
			12'hb69: tri_word = 16'h496f;
			12'hb6a: tri_word = 16'h495f;
			12'hb6b: tri_word = 16'h494f;
			12'hb6c: tri_word = 16'h493f;
			12'hb6d: tri_word = 16'h492f;
			12'hb6e: tri_word = 16'h491f;
			12'hb6f: tri_word = 16'h490f;
			12'hb70: tri_word = 16'h48ff;
			12'hb71: tri_word = 16'h48ef;
			12'hb72: tri_word = 16'h48df;
			12'hb73: tri_word = 16'h48cf;
			12'hb74: tri_word = 16'h48bf;
			12'hb75: tri_word = 16'h48af;
			12'hb76: tri_word = 16'h489f;
			12'hb77: tri_word = 16'h488f;
			12'hb78: tri_word = 16'h487f;
			12'hb79: tri_word = 16'h486f;
			12'hb7a: tri_word = 16'h485f;
			12'hb7b: tri_word = 16'h484f;
			12'hb7c: tri_word = 16'h483f;
			12'hb7d: tri_word = 16'h482f;
			12'hb7e: tri_word = 16'h481f;
			12'hb7f: tri_word = 16'h480f;
			12'hb80: tri_word = 16'h47ff;
			12'hb81: tri_word = 16'h47ef;
			12'hb82: tri_word = 16'h47df;
			12'hb83: tri_word = 16'h47cf;
			12'hb84: tri_word = 16'h47bf;
			12'hb85: tri_word = 16'h47af;
			12'hb86: tri_word = 16'h479f;
			12'hb87: tri_word = 16'h478f;
			12'hb88: tri_word = 16'h477f;
			12'hb89: tri_word = 16'h476f;
			12'hb8a: tri_word = 16'h475f;
			12'hb8b: tri_word = 16'h474f;
			12'hb8c: tri_word = 16'h473f;
			12'hb8d: tri_word = 16'h472f;
			12'hb8e: tri_word = 16'h471f;
			12'hb8f: tri_word = 16'h470f;
			12'hb90: tri_word = 16'h46ff;
			12'hb91: tri_word = 16'h46ef;
			12'hb92: tri_word = 16'h46df;
			12'hb93: tri_word = 16'h46cf;
			12'hb94: tri_word = 16'h46bf;
			12'hb95: tri_word = 16'h46af;
			12'hb96: tri_word = 16'h469f;
			12'hb97: tri_word = 16'h468f;
			12'hb98: tri_word = 16'h467f;
			12'hb99: tri_word = 16'h466f;
			12'hb9a: tri_word = 16'h465f;
			12'hb9b: tri_word = 16'h464f;
			12'hb9c: tri_word = 16'h463f;
			12'hb9d: tri_word = 16'h462f;
			12'hb9e: tri_word = 16'h461f;
			12'hb9f: tri_word = 16'h460f;
			12'hba0: tri_word = 16'h45ff;
			12'hba1: tri_word = 16'h45ef;
			12'hba2: tri_word = 16'h45df;
			12'hba3: tri_word = 16'h45cf;
			12'hba4: tri_word = 16'h45bf;
			12'hba5: tri_word = 16'h45af;
			12'hba6: tri_word = 16'h459f;
			12'hba7: tri_word = 16'h458f;
			12'hba8: tri_word = 16'h457f;
			12'hba9: tri_word = 16'h456f;
			12'hbaa: tri_word = 16'h455f;
			12'hbab: tri_word = 16'h454f;
			12'hbac: tri_word = 16'h453f;
			12'hbad: tri_word = 16'h452f;
			12'hbae: tri_word = 16'h451f;
			12'hbaf: tri_word = 16'h450f;
			12'hbb0: tri_word = 16'h44ff;
			12'hbb1: tri_word = 16'h44ef;
			12'hbb2: tri_word = 16'h44df;
			12'hbb3: tri_word = 16'h44cf;
			12'hbb4: tri_word = 16'h44bf;
			12'hbb5: tri_word = 16'h44af;
			12'hbb6: tri_word = 16'h449f;
			12'hbb7: tri_word = 16'h448f;
			12'hbb8: tri_word = 16'h447f;
			12'hbb9: tri_word = 16'h446f;
			12'hbba: tri_word = 16'h445f;
			12'hbbb: tri_word = 16'h444f;
			12'hbbc: tri_word = 16'h443f;
			12'hbbd: tri_word = 16'h442f;
			12'hbbe: tri_word = 16'h441f;
			12'hbbf: tri_word = 16'h440f;
			12'hbc0: tri_word = 16'h43ff;
			12'hbc1: tri_word = 16'h43ef;
			12'hbc2: tri_word = 16'h43df;
			12'hbc3: tri_word = 16'h43cf;
			12'hbc4: tri_word = 16'h43bf;
			12'hbc5: tri_word = 16'h43af;
			12'hbc6: tri_word = 16'h439f;
			12'hbc7: tri_word = 16'h438f;
			12'hbc8: tri_word = 16'h437f;
			12'hbc9: tri_word = 16'h436f;
			12'hbca: tri_word = 16'h435f;
			12'hbcb: tri_word = 16'h434f;
			12'hbcc: tri_word = 16'h433f;
			12'hbcd: tri_word = 16'h432f;
			12'hbce: tri_word = 16'h431f;
			12'hbcf: tri_word = 16'h430f;
			12'hbd0: tri_word = 16'h42ff;
			12'hbd1: tri_word = 16'h42ef;
			12'hbd2: tri_word = 16'h42df;
			12'hbd3: tri_word = 16'h42cf;
			12'hbd4: tri_word = 16'h42bf;
			12'hbd5: tri_word = 16'h42af;
			12'hbd6: tri_word = 16'h429f;
			12'hbd7: tri_word = 16'h428f;
			12'hbd8: tri_word = 16'h427f;
			12'hbd9: tri_word = 16'h426f;
			12'hbda: tri_word = 16'h425f;
			12'hbdb: tri_word = 16'h424f;
			12'hbdc: tri_word = 16'h423f;
			12'hbdd: tri_word = 16'h422f;
			12'hbde: tri_word = 16'h421f;
			12'hbdf: tri_word = 16'h420f;
			12'hbe0: tri_word = 16'h41ff;
			12'hbe1: tri_word = 16'h41ef;
			12'hbe2: tri_word = 16'h41df;
			12'hbe3: tri_word = 16'h41cf;
			12'hbe4: tri_word = 16'h41bf;
			12'hbe5: tri_word = 16'h41af;
			12'hbe6: tri_word = 16'h419f;
			12'hbe7: tri_word = 16'h418f;
			12'hbe8: tri_word = 16'h417f;
			12'hbe9: tri_word = 16'h416f;
			12'hbea: tri_word = 16'h415f;
			12'hbeb: tri_word = 16'h414f;
			12'hbec: tri_word = 16'h413f;
			12'hbed: tri_word = 16'h412f;
			12'hbee: tri_word = 16'h411f;
			12'hbef: tri_word = 16'h410f;
			12'hbf0: tri_word = 16'h40ff;
			12'hbf1: tri_word = 16'h40ef;
			12'hbf2: tri_word = 16'h40df;
			12'hbf3: tri_word = 16'h40cf;
			12'hbf4: tri_word = 16'h40bf;
			12'hbf5: tri_word = 16'h40af;
			12'hbf6: tri_word = 16'h409f;
			12'hbf7: tri_word = 16'h408f;
			12'hbf8: tri_word = 16'h407f;
			12'hbf9: tri_word = 16'h406f;
			12'hbfa: tri_word = 16'h405f;
			12'hbfb: tri_word = 16'h404f;
			12'hbfc: tri_word = 16'h403f;
			12'hbfd: tri_word = 16'h402f;
			12'hbfe: tri_word = 16'h401f;
			12'hbff: tri_word = 16'h400f;
			12'hc00: tri_word = 16'h3fff;
			12'hc01: tri_word = 16'h3fef;
			12'hc02: tri_word = 16'h3fdf;
			12'hc03: tri_word = 16'h3fcf;
			12'hc04: tri_word = 16'h3fbf;
			12'hc05: tri_word = 16'h3faf;
			12'hc06: tri_word = 16'h3f9f;
			12'hc07: tri_word = 16'h3f8f;
			12'hc08: tri_word = 16'h3f7f;
			12'hc09: tri_word = 16'h3f6f;
			12'hc0a: tri_word = 16'h3f5f;
			12'hc0b: tri_word = 16'h3f4f;
			12'hc0c: tri_word = 16'h3f3f;
			12'hc0d: tri_word = 16'h3f2f;
			12'hc0e: tri_word = 16'h3f1f;
			12'hc0f: tri_word = 16'h3f0f;
			12'hc10: tri_word = 16'h3eff;
			12'hc11: tri_word = 16'h3eef;
			12'hc12: tri_word = 16'h3edf;
			12'hc13: tri_word = 16'h3ecf;
			12'hc14: tri_word = 16'h3ebf;
			12'hc15: tri_word = 16'h3eaf;
			12'hc16: tri_word = 16'h3e9f;
			12'hc17: tri_word = 16'h3e8f;
			12'hc18: tri_word = 16'h3e7f;
			12'hc19: tri_word = 16'h3e6f;
			12'hc1a: tri_word = 16'h3e5f;
			12'hc1b: tri_word = 16'h3e4f;
			12'hc1c: tri_word = 16'h3e3f;
			12'hc1d: tri_word = 16'h3e2f;
			12'hc1e: tri_word = 16'h3e1f;
			12'hc1f: tri_word = 16'h3e0f;
			12'hc20: tri_word = 16'h3dff;
			12'hc21: tri_word = 16'h3def;
			12'hc22: tri_word = 16'h3ddf;
			12'hc23: tri_word = 16'h3dcf;
			12'hc24: tri_word = 16'h3dbf;
			12'hc25: tri_word = 16'h3daf;
			12'hc26: tri_word = 16'h3d9f;
			12'hc27: tri_word = 16'h3d8f;
			12'hc28: tri_word = 16'h3d7f;
			12'hc29: tri_word = 16'h3d6f;
			12'hc2a: tri_word = 16'h3d5f;
			12'hc2b: tri_word = 16'h3d4f;
			12'hc2c: tri_word = 16'h3d3f;
			12'hc2d: tri_word = 16'h3d2f;
			12'hc2e: tri_word = 16'h3d1f;
			12'hc2f: tri_word = 16'h3d0f;
			12'hc30: tri_word = 16'h3cff;
			12'hc31: tri_word = 16'h3cef;
			12'hc32: tri_word = 16'h3cdf;
			12'hc33: tri_word = 16'h3ccf;
			12'hc34: tri_word = 16'h3cbf;
			12'hc35: tri_word = 16'h3caf;
			12'hc36: tri_word = 16'h3c9f;
			12'hc37: tri_word = 16'h3c8f;
			12'hc38: tri_word = 16'h3c7f;
			12'hc39: tri_word = 16'h3c6f;
			12'hc3a: tri_word = 16'h3c5f;
			12'hc3b: tri_word = 16'h3c4f;
			12'hc3c: tri_word = 16'h3c3f;
			12'hc3d: tri_word = 16'h3c2f;
			12'hc3e: tri_word = 16'h3c1f;
			12'hc3f: tri_word = 16'h3c0f;
			12'hc40: tri_word = 16'h3bff;
			12'hc41: tri_word = 16'h3bef;
			12'hc42: tri_word = 16'h3bdf;
			12'hc43: tri_word = 16'h3bcf;
			12'hc44: tri_word = 16'h3bbf;
			12'hc45: tri_word = 16'h3baf;
			12'hc46: tri_word = 16'h3b9f;
			12'hc47: tri_word = 16'h3b8f;
			12'hc48: tri_word = 16'h3b7f;
			12'hc49: tri_word = 16'h3b6f;
			12'hc4a: tri_word = 16'h3b5f;
			12'hc4b: tri_word = 16'h3b4f;
			12'hc4c: tri_word = 16'h3b3f;
			12'hc4d: tri_word = 16'h3b2f;
			12'hc4e: tri_word = 16'h3b1f;
			12'hc4f: tri_word = 16'h3b0f;
			12'hc50: tri_word = 16'h3aff;
			12'hc51: tri_word = 16'h3aef;
			12'hc52: tri_word = 16'h3adf;
			12'hc53: tri_word = 16'h3acf;
			12'hc54: tri_word = 16'h3abf;
			12'hc55: tri_word = 16'h3aaf;
			12'hc56: tri_word = 16'h3a9f;
			12'hc57: tri_word = 16'h3a8f;
			12'hc58: tri_word = 16'h3a7f;
			12'hc59: tri_word = 16'h3a6f;
			12'hc5a: tri_word = 16'h3a5f;
			12'hc5b: tri_word = 16'h3a4f;
			12'hc5c: tri_word = 16'h3a3f;
			12'hc5d: tri_word = 16'h3a2f;
			12'hc5e: tri_word = 16'h3a1f;
			12'hc5f: tri_word = 16'h3a0f;
			12'hc60: tri_word = 16'h39ff;
			12'hc61: tri_word = 16'h39ef;
			12'hc62: tri_word = 16'h39df;
			12'hc63: tri_word = 16'h39cf;
			12'hc64: tri_word = 16'h39bf;
			12'hc65: tri_word = 16'h39af;
			12'hc66: tri_word = 16'h399f;
			12'hc67: tri_word = 16'h398f;
			12'hc68: tri_word = 16'h397f;
			12'hc69: tri_word = 16'h396f;
			12'hc6a: tri_word = 16'h395f;
			12'hc6b: tri_word = 16'h394f;
			12'hc6c: tri_word = 16'h393f;
			12'hc6d: tri_word = 16'h392f;
			12'hc6e: tri_word = 16'h391f;
			12'hc6f: tri_word = 16'h390f;
			12'hc70: tri_word = 16'h38ff;
			12'hc71: tri_word = 16'h38ef;
			12'hc72: tri_word = 16'h38df;
			12'hc73: tri_word = 16'h38cf;
			12'hc74: tri_word = 16'h38bf;
			12'hc75: tri_word = 16'h38af;
			12'hc76: tri_word = 16'h389f;
			12'hc77: tri_word = 16'h388f;
			12'hc78: tri_word = 16'h387f;
			12'hc79: tri_word = 16'h386f;
			12'hc7a: tri_word = 16'h385f;
			12'hc7b: tri_word = 16'h384f;
			12'hc7c: tri_word = 16'h383f;
			12'hc7d: tri_word = 16'h382f;
			12'hc7e: tri_word = 16'h381f;
			12'hc7f: tri_word = 16'h380f;
			12'hc80: tri_word = 16'h37ff;
			12'hc81: tri_word = 16'h37ef;
			12'hc82: tri_word = 16'h37df;
			12'hc83: tri_word = 16'h37cf;
			12'hc84: tri_word = 16'h37bf;
			12'hc85: tri_word = 16'h37af;
			12'hc86: tri_word = 16'h379f;
			12'hc87: tri_word = 16'h378f;
			12'hc88: tri_word = 16'h377f;
			12'hc89: tri_word = 16'h376f;
			12'hc8a: tri_word = 16'h375f;
			12'hc8b: tri_word = 16'h374f;
			12'hc8c: tri_word = 16'h373f;
			12'hc8d: tri_word = 16'h372f;
			12'hc8e: tri_word = 16'h371f;
			12'hc8f: tri_word = 16'h370f;
			12'hc90: tri_word = 16'h36ff;
			12'hc91: tri_word = 16'h36ef;
			12'hc92: tri_word = 16'h36df;
			12'hc93: tri_word = 16'h36cf;
			12'hc94: tri_word = 16'h36bf;
			12'hc95: tri_word = 16'h36af;
			12'hc96: tri_word = 16'h369f;
			12'hc97: tri_word = 16'h368f;
			12'hc98: tri_word = 16'h367f;
			12'hc99: tri_word = 16'h366f;
			12'hc9a: tri_word = 16'h365f;
			12'hc9b: tri_word = 16'h364f;
			12'hc9c: tri_word = 16'h363f;
			12'hc9d: tri_word = 16'h362f;
			12'hc9e: tri_word = 16'h361f;
			12'hc9f: tri_word = 16'h360f;
			12'hca0: tri_word = 16'h35ff;
			12'hca1: tri_word = 16'h35ef;
			12'hca2: tri_word = 16'h35df;
			12'hca3: tri_word = 16'h35cf;
			12'hca4: tri_word = 16'h35bf;
			12'hca5: tri_word = 16'h35af;
			12'hca6: tri_word = 16'h359f;
			12'hca7: tri_word = 16'h358f;
			12'hca8: tri_word = 16'h357f;
			12'hca9: tri_word = 16'h356f;
			12'hcaa: tri_word = 16'h355f;
			12'hcab: tri_word = 16'h354f;
			12'hcac: tri_word = 16'h353f;
			12'hcad: tri_word = 16'h352f;
			12'hcae: tri_word = 16'h351f;
			12'hcaf: tri_word = 16'h350f;
			12'hcb0: tri_word = 16'h34ff;
			12'hcb1: tri_word = 16'h34ef;
			12'hcb2: tri_word = 16'h34df;
			12'hcb3: tri_word = 16'h34cf;
			12'hcb4: tri_word = 16'h34bf;
			12'hcb5: tri_word = 16'h34af;
			12'hcb6: tri_word = 16'h349f;
			12'hcb7: tri_word = 16'h348f;
			12'hcb8: tri_word = 16'h347f;
			12'hcb9: tri_word = 16'h346f;
			12'hcba: tri_word = 16'h345f;
			12'hcbb: tri_word = 16'h344f;
			12'hcbc: tri_word = 16'h343f;
			12'hcbd: tri_word = 16'h342f;
			12'hcbe: tri_word = 16'h341f;
			12'hcbf: tri_word = 16'h340f;
			12'hcc0: tri_word = 16'h33ff;
			12'hcc1: tri_word = 16'h33ef;
			12'hcc2: tri_word = 16'h33df;
			12'hcc3: tri_word = 16'h33cf;
			12'hcc4: tri_word = 16'h33bf;
			12'hcc5: tri_word = 16'h33af;
			12'hcc6: tri_word = 16'h339f;
			12'hcc7: tri_word = 16'h338f;
			12'hcc8: tri_word = 16'h337f;
			12'hcc9: tri_word = 16'h336f;
			12'hcca: tri_word = 16'h335f;
			12'hccb: tri_word = 16'h334f;
			12'hccc: tri_word = 16'h333f;
			12'hccd: tri_word = 16'h332f;
			12'hcce: tri_word = 16'h331f;
			12'hccf: tri_word = 16'h330f;
			12'hcd0: tri_word = 16'h32ff;
			12'hcd1: tri_word = 16'h32ef;
			12'hcd2: tri_word = 16'h32df;
			12'hcd3: tri_word = 16'h32cf;
			12'hcd4: tri_word = 16'h32bf;
			12'hcd5: tri_word = 16'h32af;
			12'hcd6: tri_word = 16'h329f;
			12'hcd7: tri_word = 16'h328f;
			12'hcd8: tri_word = 16'h327f;
			12'hcd9: tri_word = 16'h326f;
			12'hcda: tri_word = 16'h325f;
			12'hcdb: tri_word = 16'h324f;
			12'hcdc: tri_word = 16'h323f;
			12'hcdd: tri_word = 16'h322f;
			12'hcde: tri_word = 16'h321f;
			12'hcdf: tri_word = 16'h320f;
			12'hce0: tri_word = 16'h31ff;
			12'hce1: tri_word = 16'h31ef;
			12'hce2: tri_word = 16'h31df;
			12'hce3: tri_word = 16'h31cf;
			12'hce4: tri_word = 16'h31bf;
			12'hce5: tri_word = 16'h31af;
			12'hce6: tri_word = 16'h319f;
			12'hce7: tri_word = 16'h318f;
			12'hce8: tri_word = 16'h317f;
			12'hce9: tri_word = 16'h316f;
			12'hcea: tri_word = 16'h315f;
			12'hceb: tri_word = 16'h314f;
			12'hcec: tri_word = 16'h313f;
			12'hced: tri_word = 16'h312f;
			12'hcee: tri_word = 16'h311f;
			12'hcef: tri_word = 16'h310f;
			12'hcf0: tri_word = 16'h30ff;
			12'hcf1: tri_word = 16'h30ef;
			12'hcf2: tri_word = 16'h30df;
			12'hcf3: tri_word = 16'h30cf;
			12'hcf4: tri_word = 16'h30bf;
			12'hcf5: tri_word = 16'h30af;
			12'hcf6: tri_word = 16'h309f;
			12'hcf7: tri_word = 16'h308f;
			12'hcf8: tri_word = 16'h307f;
			12'hcf9: tri_word = 16'h306f;
			12'hcfa: tri_word = 16'h305f;
			12'hcfb: tri_word = 16'h304f;
			12'hcfc: tri_word = 16'h303f;
			12'hcfd: tri_word = 16'h302f;
			12'hcfe: tri_word = 16'h301f;
			12'hcff: tri_word = 16'h300f;
			12'hd00: tri_word = 16'h2fff;
			12'hd01: tri_word = 16'h2fef;
			12'hd02: tri_word = 16'h2fdf;
			12'hd03: tri_word = 16'h2fcf;
			12'hd04: tri_word = 16'h2fbf;
			12'hd05: tri_word = 16'h2faf;
			12'hd06: tri_word = 16'h2f9f;
			12'hd07: tri_word = 16'h2f8f;
			12'hd08: tri_word = 16'h2f7f;
			12'hd09: tri_word = 16'h2f6f;
			12'hd0a: tri_word = 16'h2f5f;
			12'hd0b: tri_word = 16'h2f4f;
			12'hd0c: tri_word = 16'h2f3f;
			12'hd0d: tri_word = 16'h2f2f;
			12'hd0e: tri_word = 16'h2f1f;
			12'hd0f: tri_word = 16'h2f0f;
			12'hd10: tri_word = 16'h2eff;
			12'hd11: tri_word = 16'h2eef;
			12'hd12: tri_word = 16'h2edf;
			12'hd13: tri_word = 16'h2ecf;
			12'hd14: tri_word = 16'h2ebf;
			12'hd15: tri_word = 16'h2eaf;
			12'hd16: tri_word = 16'h2e9f;
			12'hd17: tri_word = 16'h2e8f;
			12'hd18: tri_word = 16'h2e7f;
			12'hd19: tri_word = 16'h2e6f;
			12'hd1a: tri_word = 16'h2e5f;
			12'hd1b: tri_word = 16'h2e4f;
			12'hd1c: tri_word = 16'h2e3f;
			12'hd1d: tri_word = 16'h2e2f;
			12'hd1e: tri_word = 16'h2e1f;
			12'hd1f: tri_word = 16'h2e0f;
			12'hd20: tri_word = 16'h2dff;
			12'hd21: tri_word = 16'h2def;
			12'hd22: tri_word = 16'h2ddf;
			12'hd23: tri_word = 16'h2dcf;
			12'hd24: tri_word = 16'h2dbf;
			12'hd25: tri_word = 16'h2daf;
			12'hd26: tri_word = 16'h2d9f;
			12'hd27: tri_word = 16'h2d8f;
			12'hd28: tri_word = 16'h2d7f;
			12'hd29: tri_word = 16'h2d6f;
			12'hd2a: tri_word = 16'h2d5f;
			12'hd2b: tri_word = 16'h2d4f;
			12'hd2c: tri_word = 16'h2d3f;
			12'hd2d: tri_word = 16'h2d2f;
			12'hd2e: tri_word = 16'h2d1f;
			12'hd2f: tri_word = 16'h2d0f;
			12'hd30: tri_word = 16'h2cff;
			12'hd31: tri_word = 16'h2cef;
			12'hd32: tri_word = 16'h2cdf;
			12'hd33: tri_word = 16'h2ccf;
			12'hd34: tri_word = 16'h2cbf;
			12'hd35: tri_word = 16'h2caf;
			12'hd36: tri_word = 16'h2c9f;
			12'hd37: tri_word = 16'h2c8f;
			12'hd38: tri_word = 16'h2c7f;
			12'hd39: tri_word = 16'h2c6f;
			12'hd3a: tri_word = 16'h2c5f;
			12'hd3b: tri_word = 16'h2c4f;
			12'hd3c: tri_word = 16'h2c3f;
			12'hd3d: tri_word = 16'h2c2f;
			12'hd3e: tri_word = 16'h2c1f;
			12'hd3f: tri_word = 16'h2c0f;
			12'hd40: tri_word = 16'h2bff;
			12'hd41: tri_word = 16'h2bef;
			12'hd42: tri_word = 16'h2bdf;
			12'hd43: tri_word = 16'h2bcf;
			12'hd44: tri_word = 16'h2bbf;
			12'hd45: tri_word = 16'h2baf;
			12'hd46: tri_word = 16'h2b9f;
			12'hd47: tri_word = 16'h2b8f;
			12'hd48: tri_word = 16'h2b7f;
			12'hd49: tri_word = 16'h2b6f;
			12'hd4a: tri_word = 16'h2b5f;
			12'hd4b: tri_word = 16'h2b4f;
			12'hd4c: tri_word = 16'h2b3f;
			12'hd4d: tri_word = 16'h2b2f;
			12'hd4e: tri_word = 16'h2b1f;
			12'hd4f: tri_word = 16'h2b0f;
			12'hd50: tri_word = 16'h2aff;
			12'hd51: tri_word = 16'h2aef;
			12'hd52: tri_word = 16'h2adf;
			12'hd53: tri_word = 16'h2acf;
			12'hd54: tri_word = 16'h2abf;
			12'hd55: tri_word = 16'h2aaf;
			12'hd56: tri_word = 16'h2a9f;
			12'hd57: tri_word = 16'h2a8f;
			12'hd58: tri_word = 16'h2a7f;
			12'hd59: tri_word = 16'h2a6f;
			12'hd5a: tri_word = 16'h2a5f;
			12'hd5b: tri_word = 16'h2a4f;
			12'hd5c: tri_word = 16'h2a3f;
			12'hd5d: tri_word = 16'h2a2f;
			12'hd5e: tri_word = 16'h2a1f;
			12'hd5f: tri_word = 16'h2a0f;
			12'hd60: tri_word = 16'h29ff;
			12'hd61: tri_word = 16'h29ef;
			12'hd62: tri_word = 16'h29df;
			12'hd63: tri_word = 16'h29cf;
			12'hd64: tri_word = 16'h29bf;
			12'hd65: tri_word = 16'h29af;
			12'hd66: tri_word = 16'h299f;
			12'hd67: tri_word = 16'h298f;
			12'hd68: tri_word = 16'h297f;
			12'hd69: tri_word = 16'h296f;
			12'hd6a: tri_word = 16'h295f;
			12'hd6b: tri_word = 16'h294f;
			12'hd6c: tri_word = 16'h293f;
			12'hd6d: tri_word = 16'h292f;
			12'hd6e: tri_word = 16'h291f;
			12'hd6f: tri_word = 16'h290f;
			12'hd70: tri_word = 16'h28ff;
			12'hd71: tri_word = 16'h28ef;
			12'hd72: tri_word = 16'h28df;
			12'hd73: tri_word = 16'h28cf;
			12'hd74: tri_word = 16'h28bf;
			12'hd75: tri_word = 16'h28af;
			12'hd76: tri_word = 16'h289f;
			12'hd77: tri_word = 16'h288f;
			12'hd78: tri_word = 16'h287f;
			12'hd79: tri_word = 16'h286f;
			12'hd7a: tri_word = 16'h285f;
			12'hd7b: tri_word = 16'h284f;
			12'hd7c: tri_word = 16'h283f;
			12'hd7d: tri_word = 16'h282f;
			12'hd7e: tri_word = 16'h281f;
			12'hd7f: tri_word = 16'h280f;
			12'hd80: tri_word = 16'h27ff;
			12'hd81: tri_word = 16'h27ef;
			12'hd82: tri_word = 16'h27df;
			12'hd83: tri_word = 16'h27cf;
			12'hd84: tri_word = 16'h27bf;
			12'hd85: tri_word = 16'h27af;
			12'hd86: tri_word = 16'h279f;
			12'hd87: tri_word = 16'h278f;
			12'hd88: tri_word = 16'h277f;
			12'hd89: tri_word = 16'h276f;
			12'hd8a: tri_word = 16'h275f;
			12'hd8b: tri_word = 16'h274f;
			12'hd8c: tri_word = 16'h273f;
			12'hd8d: tri_word = 16'h272f;
			12'hd8e: tri_word = 16'h271f;
			12'hd8f: tri_word = 16'h270f;
			12'hd90: tri_word = 16'h26ff;
			12'hd91: tri_word = 16'h26ef;
			12'hd92: tri_word = 16'h26df;
			12'hd93: tri_word = 16'h26cf;
			12'hd94: tri_word = 16'h26bf;
			12'hd95: tri_word = 16'h26af;
			12'hd96: tri_word = 16'h269f;
			12'hd97: tri_word = 16'h268f;
			12'hd98: tri_word = 16'h267f;
			12'hd99: tri_word = 16'h266f;
			12'hd9a: tri_word = 16'h265f;
			12'hd9b: tri_word = 16'h264f;
			12'hd9c: tri_word = 16'h263f;
			12'hd9d: tri_word = 16'h262f;
			12'hd9e: tri_word = 16'h261f;
			12'hd9f: tri_word = 16'h260f;
			12'hda0: tri_word = 16'h25ff;
			12'hda1: tri_word = 16'h25ef;
			12'hda2: tri_word = 16'h25df;
			12'hda3: tri_word = 16'h25cf;
			12'hda4: tri_word = 16'h25bf;
			12'hda5: tri_word = 16'h25af;
			12'hda6: tri_word = 16'h259f;
			12'hda7: tri_word = 16'h258f;
			12'hda8: tri_word = 16'h257f;
			12'hda9: tri_word = 16'h256f;
			12'hdaa: tri_word = 16'h255f;
			12'hdab: tri_word = 16'h254f;
			12'hdac: tri_word = 16'h253f;
			12'hdad: tri_word = 16'h252f;
			12'hdae: tri_word = 16'h251f;
			12'hdaf: tri_word = 16'h250f;
			12'hdb0: tri_word = 16'h24ff;
			12'hdb1: tri_word = 16'h24ef;
			12'hdb2: tri_word = 16'h24df;
			12'hdb3: tri_word = 16'h24cf;
			12'hdb4: tri_word = 16'h24bf;
			12'hdb5: tri_word = 16'h24af;
			12'hdb6: tri_word = 16'h249f;
			12'hdb7: tri_word = 16'h248f;
			12'hdb8: tri_word = 16'h247f;
			12'hdb9: tri_word = 16'h246f;
			12'hdba: tri_word = 16'h245f;
			12'hdbb: tri_word = 16'h244f;
			12'hdbc: tri_word = 16'h243f;
			12'hdbd: tri_word = 16'h242f;
			12'hdbe: tri_word = 16'h241f;
			12'hdbf: tri_word = 16'h240f;
			12'hdc0: tri_word = 16'h23ff;
			12'hdc1: tri_word = 16'h23ef;
			12'hdc2: tri_word = 16'h23df;
			12'hdc3: tri_word = 16'h23cf;
			12'hdc4: tri_word = 16'h23bf;
			12'hdc5: tri_word = 16'h23af;
			12'hdc6: tri_word = 16'h239f;
			12'hdc7: tri_word = 16'h238f;
			12'hdc8: tri_word = 16'h237f;
			12'hdc9: tri_word = 16'h236f;
			12'hdca: tri_word = 16'h235f;
			12'hdcb: tri_word = 16'h234f;
			12'hdcc: tri_word = 16'h233f;
			12'hdcd: tri_word = 16'h232f;
			12'hdce: tri_word = 16'h231f;
			12'hdcf: tri_word = 16'h230f;
			12'hdd0: tri_word = 16'h22ff;
			12'hdd1: tri_word = 16'h22ef;
			12'hdd2: tri_word = 16'h22df;
			12'hdd3: tri_word = 16'h22cf;
			12'hdd4: tri_word = 16'h22bf;
			12'hdd5: tri_word = 16'h22af;
			12'hdd6: tri_word = 16'h229f;
			12'hdd7: tri_word = 16'h228f;
			12'hdd8: tri_word = 16'h227f;
			12'hdd9: tri_word = 16'h226f;
			12'hdda: tri_word = 16'h225f;
			12'hddb: tri_word = 16'h224f;
			12'hddc: tri_word = 16'h223f;
			12'hddd: tri_word = 16'h222f;
			12'hdde: tri_word = 16'h221f;
			12'hddf: tri_word = 16'h220f;
			12'hde0: tri_word = 16'h21ff;
			12'hde1: tri_word = 16'h21ef;
			12'hde2: tri_word = 16'h21df;
			12'hde3: tri_word = 16'h21cf;
			12'hde4: tri_word = 16'h21bf;
			12'hde5: tri_word = 16'h21af;
			12'hde6: tri_word = 16'h219f;
			12'hde7: tri_word = 16'h218f;
			12'hde8: tri_word = 16'h217f;
			12'hde9: tri_word = 16'h216f;
			12'hdea: tri_word = 16'h215f;
			12'hdeb: tri_word = 16'h214f;
			12'hdec: tri_word = 16'h213f;
			12'hded: tri_word = 16'h212f;
			12'hdee: tri_word = 16'h211f;
			12'hdef: tri_word = 16'h210f;
			12'hdf0: tri_word = 16'h20ff;
			12'hdf1: tri_word = 16'h20ef;
			12'hdf2: tri_word = 16'h20df;
			12'hdf3: tri_word = 16'h20cf;
			12'hdf4: tri_word = 16'h20bf;
			12'hdf5: tri_word = 16'h20af;
			12'hdf6: tri_word = 16'h209f;
			12'hdf7: tri_word = 16'h208f;
			12'hdf8: tri_word = 16'h207f;
			12'hdf9: tri_word = 16'h206f;
			12'hdfa: tri_word = 16'h205f;
			12'hdfb: tri_word = 16'h204f;
			12'hdfc: tri_word = 16'h203f;
			12'hdfd: tri_word = 16'h202f;
			12'hdfe: tri_word = 16'h201f;
			12'hdff: tri_word = 16'h200f;
			12'he00: tri_word = 16'h1fff;
			12'he01: tri_word = 16'h1fef;
			12'he02: tri_word = 16'h1fdf;
			12'he03: tri_word = 16'h1fcf;
			12'he04: tri_word = 16'h1fbf;
			12'he05: tri_word = 16'h1faf;
			12'he06: tri_word = 16'h1f9f;
			12'he07: tri_word = 16'h1f8f;
			12'he08: tri_word = 16'h1f7f;
			12'he09: tri_word = 16'h1f6f;
			12'he0a: tri_word = 16'h1f5f;
			12'he0b: tri_word = 16'h1f4f;
			12'he0c: tri_word = 16'h1f3f;
			12'he0d: tri_word = 16'h1f2f;
			12'he0e: tri_word = 16'h1f1f;
			12'he0f: tri_word = 16'h1f0f;
			12'he10: tri_word = 16'h1eff;
			12'he11: tri_word = 16'h1eef;
			12'he12: tri_word = 16'h1edf;
			12'he13: tri_word = 16'h1ecf;
			12'he14: tri_word = 16'h1ebf;
			12'he15: tri_word = 16'h1eaf;
			12'he16: tri_word = 16'h1e9f;
			12'he17: tri_word = 16'h1e8f;
			12'he18: tri_word = 16'h1e7f;
			12'he19: tri_word = 16'h1e6f;
			12'he1a: tri_word = 16'h1e5f;
			12'he1b: tri_word = 16'h1e4f;
			12'he1c: tri_word = 16'h1e3f;
			12'he1d: tri_word = 16'h1e2f;
			12'he1e: tri_word = 16'h1e1f;
			12'he1f: tri_word = 16'h1e0f;
			12'he20: tri_word = 16'h1dff;
			12'he21: tri_word = 16'h1def;
			12'he22: tri_word = 16'h1ddf;
			12'he23: tri_word = 16'h1dcf;
			12'he24: tri_word = 16'h1dbf;
			12'he25: tri_word = 16'h1daf;
			12'he26: tri_word = 16'h1d9f;
			12'he27: tri_word = 16'h1d8f;
			12'he28: tri_word = 16'h1d7f;
			12'he29: tri_word = 16'h1d6f;
			12'he2a: tri_word = 16'h1d5f;
			12'he2b: tri_word = 16'h1d4f;
			12'he2c: tri_word = 16'h1d3f;
			12'he2d: tri_word = 16'h1d2f;
			12'he2e: tri_word = 16'h1d1f;
			12'he2f: tri_word = 16'h1d0f;
			12'he30: tri_word = 16'h1cff;
			12'he31: tri_word = 16'h1cef;
			12'he32: tri_word = 16'h1cdf;
			12'he33: tri_word = 16'h1ccf;
			12'he34: tri_word = 16'h1cbf;
			12'he35: tri_word = 16'h1caf;
			12'he36: tri_word = 16'h1c9f;
			12'he37: tri_word = 16'h1c8f;
			12'he38: tri_word = 16'h1c7f;
			12'he39: tri_word = 16'h1c6f;
			12'he3a: tri_word = 16'h1c5f;
			12'he3b: tri_word = 16'h1c4f;
			12'he3c: tri_word = 16'h1c3f;
			12'he3d: tri_word = 16'h1c2f;
			12'he3e: tri_word = 16'h1c1f;
			12'he3f: tri_word = 16'h1c0f;
			12'he40: tri_word = 16'h1bff;
			12'he41: tri_word = 16'h1bef;
			12'he42: tri_word = 16'h1bdf;
			12'he43: tri_word = 16'h1bcf;
			12'he44: tri_word = 16'h1bbf;
			12'he45: tri_word = 16'h1baf;
			12'he46: tri_word = 16'h1b9f;
			12'he47: tri_word = 16'h1b8f;
			12'he48: tri_word = 16'h1b7f;
			12'he49: tri_word = 16'h1b6f;
			12'he4a: tri_word = 16'h1b5f;
			12'he4b: tri_word = 16'h1b4f;
			12'he4c: tri_word = 16'h1b3f;
			12'he4d: tri_word = 16'h1b2f;
			12'he4e: tri_word = 16'h1b1f;
			12'he4f: tri_word = 16'h1b0f;
			12'he50: tri_word = 16'h1aff;
			12'he51: tri_word = 16'h1aef;
			12'he52: tri_word = 16'h1adf;
			12'he53: tri_word = 16'h1acf;
			12'he54: tri_word = 16'h1abf;
			12'he55: tri_word = 16'h1aaf;
			12'he56: tri_word = 16'h1a9f;
			12'he57: tri_word = 16'h1a8f;
			12'he58: tri_word = 16'h1a7f;
			12'he59: tri_word = 16'h1a6f;
			12'he5a: tri_word = 16'h1a5f;
			12'he5b: tri_word = 16'h1a4f;
			12'he5c: tri_word = 16'h1a3f;
			12'he5d: tri_word = 16'h1a2f;
			12'he5e: tri_word = 16'h1a1f;
			12'he5f: tri_word = 16'h1a0f;
			12'he60: tri_word = 16'h19ff;
			12'he61: tri_word = 16'h19ef;
			12'he62: tri_word = 16'h19df;
			12'he63: tri_word = 16'h19cf;
			12'he64: tri_word = 16'h19bf;
			12'he65: tri_word = 16'h19af;
			12'he66: tri_word = 16'h199f;
			12'he67: tri_word = 16'h198f;
			12'he68: tri_word = 16'h197f;
			12'he69: tri_word = 16'h196f;
			12'he6a: tri_word = 16'h195f;
			12'he6b: tri_word = 16'h194f;
			12'he6c: tri_word = 16'h193f;
			12'he6d: tri_word = 16'h192f;
			12'he6e: tri_word = 16'h191f;
			12'he6f: tri_word = 16'h190f;
			12'he70: tri_word = 16'h18ff;
			12'he71: tri_word = 16'h18ef;
			12'he72: tri_word = 16'h18df;
			12'he73: tri_word = 16'h18cf;
			12'he74: tri_word = 16'h18bf;
			12'he75: tri_word = 16'h18af;
			12'he76: tri_word = 16'h189f;
			12'he77: tri_word = 16'h188f;
			12'he78: tri_word = 16'h187f;
			12'he79: tri_word = 16'h186f;
			12'he7a: tri_word = 16'h185f;
			12'he7b: tri_word = 16'h184f;
			12'he7c: tri_word = 16'h183f;
			12'he7d: tri_word = 16'h182f;
			12'he7e: tri_word = 16'h181f;
			12'he7f: tri_word = 16'h180f;
			12'he80: tri_word = 16'h17ff;
			12'he81: tri_word = 16'h17ef;
			12'he82: tri_word = 16'h17df;
			12'he83: tri_word = 16'h17cf;
			12'he84: tri_word = 16'h17bf;
			12'he85: tri_word = 16'h17af;
			12'he86: tri_word = 16'h179f;
			12'he87: tri_word = 16'h178f;
			12'he88: tri_word = 16'h177f;
			12'he89: tri_word = 16'h176f;
			12'he8a: tri_word = 16'h175f;
			12'he8b: tri_word = 16'h174f;
			12'he8c: tri_word = 16'h173f;
			12'he8d: tri_word = 16'h172f;
			12'he8e: tri_word = 16'h171f;
			12'he8f: tri_word = 16'h170f;
			12'he90: tri_word = 16'h16ff;
			12'he91: tri_word = 16'h16ef;
			12'he92: tri_word = 16'h16df;
			12'he93: tri_word = 16'h16cf;
			12'he94: tri_word = 16'h16bf;
			12'he95: tri_word = 16'h16af;
			12'he96: tri_word = 16'h169f;
			12'he97: tri_word = 16'h168f;
			12'he98: tri_word = 16'h167f;
			12'he99: tri_word = 16'h166f;
			12'he9a: tri_word = 16'h165f;
			12'he9b: tri_word = 16'h164f;
			12'he9c: tri_word = 16'h163f;
			12'he9d: tri_word = 16'h162f;
			12'he9e: tri_word = 16'h161f;
			12'he9f: tri_word = 16'h160f;
			12'hea0: tri_word = 16'h15ff;
			12'hea1: tri_word = 16'h15ef;
			12'hea2: tri_word = 16'h15df;
			12'hea3: tri_word = 16'h15cf;
			12'hea4: tri_word = 16'h15bf;
			12'hea5: tri_word = 16'h15af;
			12'hea6: tri_word = 16'h159f;
			12'hea7: tri_word = 16'h158f;
			12'hea8: tri_word = 16'h157f;
			12'hea9: tri_word = 16'h156f;
			12'heaa: tri_word = 16'h155f;
			12'heab: tri_word = 16'h154f;
			12'heac: tri_word = 16'h153f;
			12'head: tri_word = 16'h152f;
			12'heae: tri_word = 16'h151f;
			12'heaf: tri_word = 16'h150f;
			12'heb0: tri_word = 16'h14ff;
			12'heb1: tri_word = 16'h14ef;
			12'heb2: tri_word = 16'h14df;
			12'heb3: tri_word = 16'h14cf;
			12'heb4: tri_word = 16'h14bf;
			12'heb5: tri_word = 16'h14af;
			12'heb6: tri_word = 16'h149f;
			12'heb7: tri_word = 16'h148f;
			12'heb8: tri_word = 16'h147f;
			12'heb9: tri_word = 16'h146f;
			12'heba: tri_word = 16'h145f;
			12'hebb: tri_word = 16'h144f;
			12'hebc: tri_word = 16'h143f;
			12'hebd: tri_word = 16'h142f;
			12'hebe: tri_word = 16'h141f;
			12'hebf: tri_word = 16'h140f;
			12'hec0: tri_word = 16'h13ff;
			12'hec1: tri_word = 16'h13ef;
			12'hec2: tri_word = 16'h13df;
			12'hec3: tri_word = 16'h13cf;
			12'hec4: tri_word = 16'h13bf;
			12'hec5: tri_word = 16'h13af;
			12'hec6: tri_word = 16'h139f;
			12'hec7: tri_word = 16'h138f;
			12'hec8: tri_word = 16'h137f;
			12'hec9: tri_word = 16'h136f;
			12'heca: tri_word = 16'h135f;
			12'hecb: tri_word = 16'h134f;
			12'hecc: tri_word = 16'h133f;
			12'hecd: tri_word = 16'h132f;
			12'hece: tri_word = 16'h131f;
			12'hecf: tri_word = 16'h130f;
			12'hed0: tri_word = 16'h12ff;
			12'hed1: tri_word = 16'h12ef;
			12'hed2: tri_word = 16'h12df;
			12'hed3: tri_word = 16'h12cf;
			12'hed4: tri_word = 16'h12bf;
			12'hed5: tri_word = 16'h12af;
			12'hed6: tri_word = 16'h129f;
			12'hed7: tri_word = 16'h128f;
			12'hed8: tri_word = 16'h127f;
			12'hed9: tri_word = 16'h126f;
			12'heda: tri_word = 16'h125f;
			12'hedb: tri_word = 16'h124f;
			12'hedc: tri_word = 16'h123f;
			12'hedd: tri_word = 16'h122f;
			12'hede: tri_word = 16'h121f;
			12'hedf: tri_word = 16'h120f;
			12'hee0: tri_word = 16'h11ff;
			12'hee1: tri_word = 16'h11ef;
			12'hee2: tri_word = 16'h11df;
			12'hee3: tri_word = 16'h11cf;
			12'hee4: tri_word = 16'h11bf;
			12'hee5: tri_word = 16'h11af;
			12'hee6: tri_word = 16'h119f;
			12'hee7: tri_word = 16'h118f;
			12'hee8: tri_word = 16'h117f;
			12'hee9: tri_word = 16'h116f;
			12'heea: tri_word = 16'h115f;
			12'heeb: tri_word = 16'h114f;
			12'heec: tri_word = 16'h113f;
			12'heed: tri_word = 16'h112f;
			12'heee: tri_word = 16'h111f;
			12'heef: tri_word = 16'h110f;
			12'hef0: tri_word = 16'h10ff;
			12'hef1: tri_word = 16'h10ef;
			12'hef2: tri_word = 16'h10df;
			12'hef3: tri_word = 16'h10cf;
			12'hef4: tri_word = 16'h10bf;
			12'hef5: tri_word = 16'h10af;
			12'hef6: tri_word = 16'h109f;
			12'hef7: tri_word = 16'h108f;
			12'hef8: tri_word = 16'h107f;
			12'hef9: tri_word = 16'h106f;
			12'hefa: tri_word = 16'h105f;
			12'hefb: tri_word = 16'h104f;
			12'hefc: tri_word = 16'h103f;
			12'hefd: tri_word = 16'h102f;
			12'hefe: tri_word = 16'h101f;
			12'heff: tri_word = 16'h100f;
			12'hf00: tri_word = 16'h0fff;
			12'hf01: tri_word = 16'h0fef;
			12'hf02: tri_word = 16'h0fdf;
			12'hf03: tri_word = 16'h0fcf;
			12'hf04: tri_word = 16'h0fbf;
			12'hf05: tri_word = 16'h0faf;
			12'hf06: tri_word = 16'h0f9f;
			12'hf07: tri_word = 16'h0f8f;
			12'hf08: tri_word = 16'h0f7f;
			12'hf09: tri_word = 16'h0f6f;
			12'hf0a: tri_word = 16'h0f5f;
			12'hf0b: tri_word = 16'h0f4f;
			12'hf0c: tri_word = 16'h0f3f;
			12'hf0d: tri_word = 16'h0f2f;
			12'hf0e: tri_word = 16'h0f1f;
			12'hf0f: tri_word = 16'h0f0f;
			12'hf10: tri_word = 16'h0eff;
			12'hf11: tri_word = 16'h0eef;
			12'hf12: tri_word = 16'h0edf;
			12'hf13: tri_word = 16'h0ecf;
			12'hf14: tri_word = 16'h0ebf;
			12'hf15: tri_word = 16'h0eaf;
			12'hf16: tri_word = 16'h0e9f;
			12'hf17: tri_word = 16'h0e8f;
			12'hf18: tri_word = 16'h0e7f;
			12'hf19: tri_word = 16'h0e6f;
			12'hf1a: tri_word = 16'h0e5f;
			12'hf1b: tri_word = 16'h0e4f;
			12'hf1c: tri_word = 16'h0e3f;
			12'hf1d: tri_word = 16'h0e2f;
			12'hf1e: tri_word = 16'h0e1f;
			12'hf1f: tri_word = 16'h0e0f;
			12'hf20: tri_word = 16'h0dff;
			12'hf21: tri_word = 16'h0def;
			12'hf22: tri_word = 16'h0ddf;
			12'hf23: tri_word = 16'h0dcf;
			12'hf24: tri_word = 16'h0dbf;
			12'hf25: tri_word = 16'h0daf;
			12'hf26: tri_word = 16'h0d9f;
			12'hf27: tri_word = 16'h0d8f;
			12'hf28: tri_word = 16'h0d7f;
			12'hf29: tri_word = 16'h0d6f;
			12'hf2a: tri_word = 16'h0d5f;
			12'hf2b: tri_word = 16'h0d4f;
			12'hf2c: tri_word = 16'h0d3f;
			12'hf2d: tri_word = 16'h0d2f;
			12'hf2e: tri_word = 16'h0d1f;
			12'hf2f: tri_word = 16'h0d0f;
			12'hf30: tri_word = 16'h0cff;
			12'hf31: tri_word = 16'h0cef;
			12'hf32: tri_word = 16'h0cdf;
			12'hf33: tri_word = 16'h0ccf;
			12'hf34: tri_word = 16'h0cbf;
			12'hf35: tri_word = 16'h0caf;
			12'hf36: tri_word = 16'h0c9f;
			12'hf37: tri_word = 16'h0c8f;
			12'hf38: tri_word = 16'h0c7f;
			12'hf39: tri_word = 16'h0c6f;
			12'hf3a: tri_word = 16'h0c5f;
			12'hf3b: tri_word = 16'h0c4f;
			12'hf3c: tri_word = 16'h0c3f;
			12'hf3d: tri_word = 16'h0c2f;
			12'hf3e: tri_word = 16'h0c1f;
			12'hf3f: tri_word = 16'h0c0f;
			12'hf40: tri_word = 16'h0bff;
			12'hf41: tri_word = 16'h0bef;
			12'hf42: tri_word = 16'h0bdf;
			12'hf43: tri_word = 16'h0bcf;
			12'hf44: tri_word = 16'h0bbf;
			12'hf45: tri_word = 16'h0baf;
			12'hf46: tri_word = 16'h0b9f;
			12'hf47: tri_word = 16'h0b8f;
			12'hf48: tri_word = 16'h0b7f;
			12'hf49: tri_word = 16'h0b6f;
			12'hf4a: tri_word = 16'h0b5f;
			12'hf4b: tri_word = 16'h0b4f;
			12'hf4c: tri_word = 16'h0b3f;
			12'hf4d: tri_word = 16'h0b2f;
			12'hf4e: tri_word = 16'h0b1f;
			12'hf4f: tri_word = 16'h0b0f;
			12'hf50: tri_word = 16'h0aff;
			12'hf51: tri_word = 16'h0aef;
			12'hf52: tri_word = 16'h0adf;
			12'hf53: tri_word = 16'h0acf;
			12'hf54: tri_word = 16'h0abf;
			12'hf55: tri_word = 16'h0aaf;
			12'hf56: tri_word = 16'h0a9f;
			12'hf57: tri_word = 16'h0a8f;
			12'hf58: tri_word = 16'h0a7f;
			12'hf59: tri_word = 16'h0a6f;
			12'hf5a: tri_word = 16'h0a5f;
			12'hf5b: tri_word = 16'h0a4f;
			12'hf5c: tri_word = 16'h0a3f;
			12'hf5d: tri_word = 16'h0a2f;
			12'hf5e: tri_word = 16'h0a1f;
			12'hf5f: tri_word = 16'h0a0f;
			12'hf60: tri_word = 16'h09ff;
			12'hf61: tri_word = 16'h09ef;
			12'hf62: tri_word = 16'h09df;
			12'hf63: tri_word = 16'h09cf;
			12'hf64: tri_word = 16'h09bf;
			12'hf65: tri_word = 16'h09af;
			12'hf66: tri_word = 16'h099f;
			12'hf67: tri_word = 16'h098f;
			12'hf68: tri_word = 16'h097f;
			12'hf69: tri_word = 16'h096f;
			12'hf6a: tri_word = 16'h095f;
			12'hf6b: tri_word = 16'h094f;
			12'hf6c: tri_word = 16'h093f;
			12'hf6d: tri_word = 16'h092f;
			12'hf6e: tri_word = 16'h091f;
			12'hf6f: tri_word = 16'h090f;
			12'hf70: tri_word = 16'h08ff;
			12'hf71: tri_word = 16'h08ef;
			12'hf72: tri_word = 16'h08df;
			12'hf73: tri_word = 16'h08cf;
			12'hf74: tri_word = 16'h08bf;
			12'hf75: tri_word = 16'h08af;
			12'hf76: tri_word = 16'h089f;
			12'hf77: tri_word = 16'h088f;
			12'hf78: tri_word = 16'h087f;
			12'hf79: tri_word = 16'h086f;
			12'hf7a: tri_word = 16'h085f;
			12'hf7b: tri_word = 16'h084f;
			12'hf7c: tri_word = 16'h083f;
			12'hf7d: tri_word = 16'h082f;
			12'hf7e: tri_word = 16'h081f;
			12'hf7f: tri_word = 16'h080f;
			12'hf80: tri_word = 16'h07ff;
			12'hf81: tri_word = 16'h07ef;
			12'hf82: tri_word = 16'h07df;
			12'hf83: tri_word = 16'h07cf;
			12'hf84: tri_word = 16'h07bf;
			12'hf85: tri_word = 16'h07af;
			12'hf86: tri_word = 16'h079f;
			12'hf87: tri_word = 16'h078f;
			12'hf88: tri_word = 16'h077f;
			12'hf89: tri_word = 16'h076f;
			12'hf8a: tri_word = 16'h075f;
			12'hf8b: tri_word = 16'h074f;
			12'hf8c: tri_word = 16'h073f;
			12'hf8d: tri_word = 16'h072f;
			12'hf8e: tri_word = 16'h071f;
			12'hf8f: tri_word = 16'h070f;
			12'hf90: tri_word = 16'h06ff;
			12'hf91: tri_word = 16'h06ef;
			12'hf92: tri_word = 16'h06df;
			12'hf93: tri_word = 16'h06cf;
			12'hf94: tri_word = 16'h06bf;
			12'hf95: tri_word = 16'h06af;
			12'hf96: tri_word = 16'h069f;
			12'hf97: tri_word = 16'h068f;
			12'hf98: tri_word = 16'h067f;
			12'hf99: tri_word = 16'h066f;
			12'hf9a: tri_word = 16'h065f;
			12'hf9b: tri_word = 16'h064f;
			12'hf9c: tri_word = 16'h063f;
			12'hf9d: tri_word = 16'h062f;
			12'hf9e: tri_word = 16'h061f;
			12'hf9f: tri_word = 16'h060f;
			12'hfa0: tri_word = 16'h05ff;
			12'hfa1: tri_word = 16'h05ef;
			12'hfa2: tri_word = 16'h05df;
			12'hfa3: tri_word = 16'h05cf;
			12'hfa4: tri_word = 16'h05bf;
			12'hfa5: tri_word = 16'h05af;
			12'hfa6: tri_word = 16'h059f;
			12'hfa7: tri_word = 16'h058f;
			12'hfa8: tri_word = 16'h057f;
			12'hfa9: tri_word = 16'h056f;
			12'hfaa: tri_word = 16'h055f;
			12'hfab: tri_word = 16'h054f;
			12'hfac: tri_word = 16'h053f;
			12'hfad: tri_word = 16'h052f;
			12'hfae: tri_word = 16'h051f;
			12'hfaf: tri_word = 16'h050f;
			12'hfb0: tri_word = 16'h04ff;
			12'hfb1: tri_word = 16'h04ef;
			12'hfb2: tri_word = 16'h04df;
			12'hfb3: tri_word = 16'h04cf;
			12'hfb4: tri_word = 16'h04bf;
			12'hfb5: tri_word = 16'h04af;
			12'hfb6: tri_word = 16'h049f;
			12'hfb7: tri_word = 16'h048f;
			12'hfb8: tri_word = 16'h047f;
			12'hfb9: tri_word = 16'h046f;
			12'hfba: tri_word = 16'h045f;
			12'hfbb: tri_word = 16'h044f;
			12'hfbc: tri_word = 16'h043f;
			12'hfbd: tri_word = 16'h042f;
			12'hfbe: tri_word = 16'h041f;
			12'hfbf: tri_word = 16'h040f;
			12'hfc0: tri_word = 16'h03ff;
			12'hfc1: tri_word = 16'h03ef;
			12'hfc2: tri_word = 16'h03df;
			12'hfc3: tri_word = 16'h03cf;
			12'hfc4: tri_word = 16'h03bf;
			12'hfc5: tri_word = 16'h03af;
			12'hfc6: tri_word = 16'h039f;
			12'hfc7: tri_word = 16'h038f;
			12'hfc8: tri_word = 16'h037f;
			12'hfc9: tri_word = 16'h036f;
			12'hfca: tri_word = 16'h035f;
			12'hfcb: tri_word = 16'h034f;
			12'hfcc: tri_word = 16'h033f;
			12'hfcd: tri_word = 16'h032f;
			12'hfce: tri_word = 16'h031f;
			12'hfcf: tri_word = 16'h030f;
			12'hfd0: tri_word = 16'h02ff;
			12'hfd1: tri_word = 16'h02ef;
			12'hfd2: tri_word = 16'h02df;
			12'hfd3: tri_word = 16'h02cf;
			12'hfd4: tri_word = 16'h02bf;
			12'hfd5: tri_word = 16'h02af;
			12'hfd6: tri_word = 16'h029f;
			12'hfd7: tri_word = 16'h028f;
			12'hfd8: tri_word = 16'h027f;
			12'hfd9: tri_word = 16'h026f;
			12'hfda: tri_word = 16'h025f;
			12'hfdb: tri_word = 16'h024f;
			12'hfdc: tri_word = 16'h023f;
			12'hfdd: tri_word = 16'h022f;
			12'hfde: tri_word = 16'h021f;
			12'hfdf: tri_word = 16'h020f;
			12'hfe0: tri_word = 16'h01ff;
			12'hfe1: tri_word = 16'h01ef;
			12'hfe2: tri_word = 16'h01df;
			12'hfe3: tri_word = 16'h01cf;
			12'hfe4: tri_word = 16'h01bf;
			12'hfe5: tri_word = 16'h01af;
			12'hfe6: tri_word = 16'h019f;
			12'hfe7: tri_word = 16'h018f;
			12'hfe8: tri_word = 16'h017f;
			12'hfe9: tri_word = 16'h016f;
			12'hfea: tri_word = 16'h015f;
			12'hfeb: tri_word = 16'h014f;
			12'hfec: tri_word = 16'h013f;
			12'hfed: tri_word = 16'h012f;
			12'hfee: tri_word = 16'h011f;
			12'hfef: tri_word = 16'h010f;
			12'hff0: tri_word = 16'h00ff;
			12'hff1: tri_word = 16'h00ef;
			12'hff2: tri_word = 16'h00df;
			12'hff3: tri_word = 16'h00cf;
			12'hff4: tri_word = 16'h00bf;
			12'hff5: tri_word = 16'h00af;
			12'hff6: tri_word = 16'h009f;
			12'hff7: tri_word = 16'h008f;
			12'hff8: tri_word = 16'h007f;
			12'hff9: tri_word = 16'h006f;
			12'hffa: tri_word = 16'h005f;
			12'hffb: tri_word = 16'h004f;
			12'hffc: tri_word = 16'h003f;
			12'hffd: tri_word = 16'h002f;
			12'hffe: tri_word = 16'h001f;
			12'hfff: tri_word = 16'h000f;
			default: tri_word = 16'h0000;
		endcase 
	end
endmodule